`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Montek Singh
// 10/22/2020
//
// PLEASE README!
// ==============
//
// This is a self-checking tester for your full MIPS processor 
// plus VGA display.
//
// Use this tester carefully!  The names of your top-level input/output
// and internal signals may be different, so modify all of signal names on the
// right-hand-side of the "wire" assigments appearing above the uut
// instantiation.  Observe that the uut itself only has clock and reset inputs
// now, and no debug outputs.  Also, the parameters specifying the names of the
// memory initialization files must match the actual file names.
//
// If you decide not to use some of these internal signals for debugging, you
// may comment the relevant lines out.  Be sure to comment out the
// corresponding "ERROR_*" lines below as well.
//
// Finally, note that in my bitmap memory, each 12-bit color is encoded as
// RRRRGGGGBBBB (i.e., red is most significant).  If you have chosen a different
// order for the red/green/blue color values, you may see ERROR signals for the
// colors light up.
//
//////////////////////////////////////////////////////////////////////////////////


module project_screentest;

    // Parameters
    localparam Nchars = 4;
    localparam charcode_size = $clog2(Nchars);
    localparam bmem_size = Nchars * 256;
     
    // Inputs
    logic clk;
    logic reset;

    // Signals inside top-level module uut
    wire [31:0] pc             =uut.pc;                    // PC
    wire [31:0] instr          =uut.instr;                 // instr coming out of instr mem
    wire [31:0] mem_addr       =uut.mem_addr;              // addr sent to data mem
    wire        mem_wr         =uut.mem_wr;                // write enable for data mem
    wire [31:0] mem_readdata   =uut.mem_readdata;          // data read from data mem
    wire [31:0] mem_writedata  =uut.mem_writedata;         // write data for data mem
    wire [31:0] period         =uut.period;                // period for sound module
    wire [15:0] LED            =uut.LED;                   // light pattern for LEDs
    
    // Signals inside module uut.mips
    wire        werf           =uut.mips.werf;              // WERF = write enable for register file
    wire  [4:0] alufn          =uut.mips.alufn;             // ALU function
    wire        Z              =uut.mips.Z;                 // Zero flag

    // Signals inside module uut.mips.dp (datapath)
    wire [31:0] ReadData1      =uut.mips.dp.ReadData1;       // Reg[rs]
    wire [31:0] ReadData2      =uut.mips.dp.ReadData2;       // Reg[rt]
    wire [31:0] alu_result     =uut.mips.dp.alu_result;      // ALU's output
    wire [4:0]  reg_writeaddr  =uut.mips.dp.reg_writeaddr;   // destination register
    wire [31:0] reg_writedata  =uut.mips.dp.reg_writedata;   // write data for register file
    wire [31:0] signImm        =uut.mips.dp.signImm;         // sign-/zero-extended immediate
    wire [31:0] aluA           =uut.mips.dp.aluA;            // operand A for ALU
    wire [31:0] aluB           =uut.mips.dp.aluB;            // operand B for ALU

    // Signals inside module uut.mips.c (controller)
    wire [1:0] pcsel           =uut.mips.c.pcsel;
    wire [1:0] wasel           =uut.mips.c.wasel;
    wire sgnext                  =uut.mips.c.sgnext;
    wire bsel                  =uut.mips.c.bsel;
    wire [1:0] wdsel           =uut.mips.c.wdsel;
    wire wr                    =uut.mips.c.wr;
    wire [1:0] asel            =uut.mips.c.asel;

    // Signals related to module memIO (memory + memory-mapped IO)
    wire [10:0] smem_addr      =uut.smem_addr;             // address from vgadisplaydriver to access screen mem
    wire [charcode_size-1:0]  charcode       =uut.charcode;              // character code returned by screen mem
    wire cpu_wr                =uut.memIO.cpu_wr;
    wire dmem_wr               =uut.memIO.dmem_wr;
    wire smem_wr               =uut.memIO.smem_wr;
    wire sound_wr              =uut.memIO.sound_wr;
    wire lights_wr             =uut.memIO.lights_wr;
    wire [31:0] smem_readdata  =uut.memIO.smem_readdata;
    wire [31:0] dmem_readdata  =uut.memIO.dmem_readdata;
    wire [31:0] keyb_char      =uut.memIO.keyb_char;
    wire [31:0] accel_val      =uut.memIO.accel_val;
    wire [31:0] cpu_addr       =uut.memIO.cpu_addr;
    wire [31:0] cpu_readdata   =uut.memIO.cpu_readdata;
    wire [31:0] cpu_writedata  =uut.memIO.cpu_writedata;
    

    // Signals related to module vgadisplaydriver (display driver)
    wire hsync                 =uut.hsync;
    wire vsync                 =uut.vsync;
    wire [3:0] red             =uut.red;
    wire [3:0] green           =uut.green;
    wire [3:0] blue            =uut.blue;
    wire [9:0] x               =uut.myDisplay.x;
    wire [9:0] y               =uut.myDisplay.y;
    wire [$clog2(bmem_size)-1:0] bmem_addr      =uut.myDisplay.BitmapAddr;
    wire [11:0] bmem_color     =uut.myDisplay.RGB;
    

    // Instantiate the Unit Under Test (UUT)
    top #(
      .Nchars(Nchars),                    // number of characters/sprites
      .imem_size(1024),                   // imem size, must be >= # instructions in program
      .imem_init("imem_screentest_nopause.mem"),    // program code
      .dmem_size(1024),                   // dmem size, must be >= # words in .data of program + size of stack
      .dmem_init("dmem_test.mem")         // program data + stack space
    ) uut(
      .clk(clk), 
      .reset(reset)
    );

//
// CHECK ALL VALUES ABOVE THIS LINE
// YOU SHOULD NOT NEED TO MODIFY ANYTHING BELOW
//

    initial begin
        // Initialize Inputs
        clk = 0;
        reset = 0;
   end

   initial begin
      #0.5 clk = 0;
      forever
         #0.5 clk = ~clk;
   end
   
   initial begin
      #1000 $finish;
   end
   
   
   
   // SELF-CHECKING CODE
   
   selfcheck_nopause c();

    wire [31:0] c_pc=c.pc;
    wire [31:0] c_instr=c.instr;
    wire [31:0] c_mem_addr=c.mem_addr;
    wire        c_mem_wr=c.mem_wr;
    wire [31:0] c_mem_readdata=c.mem_readdata;
    wire [31:0] c_mem_writedata=c.mem_writedata;
    wire [31:0] c_period=c.period;
    wire [15:0] c_LED=c.LED;
    wire        c_werf=c.werf;
    wire  [4:0] c_alufn=c.alufn;
    wire        c_Z=c.Z;
    wire [31:0] c_ReadData1=c.ReadData1;
    wire [31:0] c_ReadData2=c.ReadData2;
    wire [31:0] c_alu_result=c.alu_result;
    wire [4:0]  c_reg_writeaddr=c.reg_writeaddr;
    wire [31:0] c_reg_writedata=c.reg_writedata;
    wire [31:0] c_signImm=c.signImm;
    wire [31:0] c_aluA=c.aluA;
    wire [31:0] c_aluB=c.aluB;
    wire [1:0]  c_pcsel=c.pcsel;
    wire [1:0]  c_wasel=c.wasel;
    wire        c_sgnext=c.sgnext;
    wire        c_bsel=c.bsel;
    wire [1:0]  c_wdsel=c.wdsel;
    wire        c_wr=c.wr;
    wire [1:0]  c_asel=c.asel;
    wire [10:0] c_smem_addr=c.smem_addr;
    wire [3:0]  c_charcode=c.charcode;
    wire        c_dmem_wr=c.dmem_wr;
    wire        c_smem_wr=c.smem_wr;
    wire        c_hsync=c.hsync;
    wire        c_vsync=c.vsync;
    wire [3:0]  c_red=c.red;
    wire [3:0]  c_green=c.green;
    wire [3:0]  c_blue=c.blue;
    wire [9:0]  c_x=c.x;
    wire [9:0]  c_y=c.y;
    wire [11:0] c_bmem_addr=c.bmem_addr;
    wire [11:0] c_bmem_color=c.bmem_color;
    wire c_sound_wr=c.sound_wr;
    wire c_lights_wr=c.lights_wr;
    wire [31:0] c_smem_readdata=c.smem_readdata;
    wire [31:0] c_dmem_readdata=c.dmem_readdata;
    wire [31:0] c_keyb_char=c.keyb_char;
    wire [31:0] c_accel_val=c.accel_val;
    wire [31:0] c_cpu_addr=c.cpu_addr;
    wire [31:0] c_cpu_readdata=c.cpu_readdata;
    wire [31:0] c_cpu_writedata=c.cpu_writedata;
  

  
    function mismatch;  // some trickery needed to match two values with don't cares
        input p, q;      // mismatch in a bit position is ignored if q has an 'x' in that bit
        integer p, q;
        mismatch = (((p ^ q) ^ q) !== q);
    endfunction

    wire ERROR;
    wire ERROR_pc             = mismatch(pc, c.pc) ? 1'bx : 1'b0;
    wire ERROR_instr          = mismatch(instr, c.instr) ? 1'bx : 1'b0;
    wire ERROR_mem_addr       = mismatch(mem_addr, c.mem_addr) ? 1'bx : 1'b0;
    wire ERROR_mem_wr         = mismatch(mem_wr, c.mem_wr) ? 1'bx : 1'b0;
    wire ERROR_mem_readdata   = mismatch(mem_readdata, c.mem_readdata) ? 1'bx : 1'b0;
    wire ERROR_mem_writedata  = c.mem_wr & (mismatch(mem_writedata, c.mem_writedata) ? 1'bx : 1'b0);
    wire ERROR_period         = mismatch(period, c.period) ? 1'bx : 1'b0;
    wire ERROR_LED            = mismatch(LED, c.LED) ? 1'bx : 1'b0;
    wire ERROR_werf           = mismatch(werf, c.werf) ? 1'bx : 1'b0;
    wire ERROR_alufn          = mismatch(alufn, c.alufn) ? 1'bx : 1'b0;
    wire ERROR_Z              = mismatch(Z, c.Z) ? 1'bx : 1'b0;
    wire ERROR_ReadData1      = mismatch(ReadData1, c.ReadData1) ? 1'bx : 1'b0;
    wire ERROR_ReadData2      = mismatch(ReadData2, c.ReadData2) ? 1'bx : 1'b0;
    wire ERROR_alu_result     = mismatch(alu_result, c.alu_result) ? 1'bx : 1'b0;
    wire ERROR_reg_writeaddr  = c.werf & (mismatch(reg_writeaddr, c.reg_writeaddr) ? 1'bx : 1'b0);
    wire ERROR_reg_writedata  = c.werf & (mismatch(reg_writedata, c.reg_writedata) ? 1'bx : 1'b0);
    wire ERROR_signImm        = mismatch(signImm, c.signImm) ? 1'bx : 1'b0;
    wire ERROR_aluA           = mismatch(aluA, c.aluA) ? 1'bx : 1'b0;
    wire ERROR_aluB           = mismatch(aluB, c.aluB) ? 1'bx : 1'b0;
    wire ERROR_pcsel          = mismatch(pcsel, c.pcsel) ? 1'bx : 1'b0;
    wire ERROR_wasel          = c.werf & (mismatch(wasel, c.wasel) ? 1'bx : 1'b0);
    wire ERROR_sgnext         = mismatch(sgnext, c.sgnext) ? 1'bx : 1'b0;
    wire ERROR_bsel           = mismatch(bsel, c.bsel) ? 1'bx : 1'b0;
    wire ERROR_wdsel          = mismatch(wdsel, c.wdsel) ? 1'bx : 1'b0;
    wire ERROR_wr             = mismatch(wr, c.wr) ? 1'bx : 1'b0;
    wire ERROR_asel           = mismatch(asel, c.asel) ? 1'bx : 1'b0;
    wire ERROR_smem_addr      = mismatch(smem_addr, c.smem_addr) ? 1'bx : 1'b0;
    wire ERROR_charcode       = mismatch(charcode, c.charcode) ? 1'bx : 1'b0;
    wire ERROR_dmem_wr        = mismatch(dmem_wr, c.dmem_wr) ? 1'bx : 1'b0;
    wire ERROR_smem_wr        = mismatch(smem_wr, c.smem_wr) ? 1'bx : 1'b0;
    wire ERROR_sound_wr       = mismatch(sound_wr, c.sound_wr) ? 1'bx : 1'b0;
    wire ERROR_lights_wr      = mismatch(lights_wr, c.lights_wr) ? 1'bx : 1'b0;
    wire ERROR_smem_readdata  = mismatch(smem_readdata, c.smem_readdata) ? 1'bx : 1'b0;
    wire ERROR_dmem_readdata  = mismatch(dmem_readdata, c.dmem_readdata) ? 1'bx : 1'b0;
    wire ERROR_keyb_char      = mismatch(keyb_char, c.keyb_char) ? 1'bx : 1'b0;
    wire ERROR_accel_val      = mismatch(accel_val, c.accel_val) ? 1'bx : 1'b0;
    wire ERROR_cpu_addr       = mismatch(cpu_addr, c.cpu_addr) ? 1'bx : 1'b0;
    wire ERROR_cpu_readdata   = mismatch(cpu_readdata, c.cpu_readdata) ? 1'bx : 1'b0;
    wire ERROR_cpu_writedata  = mismatch(cpu_writedata, c.cpu_writedata) ? 1'bx : 1'b0;  
    wire ERROR_hsync          = mismatch(hsync, c.hsync) ? 1'bx : 1'b0;
    wire ERROR_vsync          = mismatch(vsync, c.vsync) ? 1'bx : 1'b0;
    wire ERROR_red            = mismatch(red, c.red) ? 1'bx : 1'b0;
    wire ERROR_green          = mismatch(green, c.green) ? 1'bx : 1'b0;
    wire ERROR_blue           = mismatch(blue, c.blue) ? 1'bx : 1'b0;
    wire ERROR_x              = mismatch(x, c.x) ? 1'bx : 1'b0;
    wire ERROR_y              = mismatch(y, c.y) ? 1'bx : 1'b0;
    wire ERROR_bmem_addr      = mismatch(bmem_addr, c.bmem_addr) ? 1'bx : 1'b0;
    wire ERROR_bmem_color     = mismatch(bmem_color, c.bmem_color) ? 1'bx : 1'b0;

    assign ERROR = ERROR_pc | ERROR_instr | ERROR_mem_addr | ERROR_mem_wr | ERROR_mem_readdata 
              | ERROR_mem_writedata | ERROR_period | ERROR_LED | ERROR_werf | ERROR_alufn | ERROR_Z
              | ERROR_ReadData1 | ERROR_ReadData2 | ERROR_alu_result | ERROR_reg_writeaddr
              | ERROR_reg_writedata | ERROR_signImm | ERROR_aluA | ERROR_aluB
              | ERROR_pcsel | ERROR_wasel | ERROR_sgnext | ERROR_bsel | ERROR_wdsel | ERROR_wr | ERROR_asel
              | ERROR_smem_addr | ERROR_charcode | ERROR_dmem_wr | ERROR_smem_wr 
              | ERROR_sound_wr | ERROR_lights_wr | ERROR_smem_readdata | ERROR_dmem_readdata
              | ERROR_keyb_char | ERROR_accel_val | ERROR_cpu_addr | ERROR_cpu_readdata | ERROR_cpu_writedata
              | ERROR_hsync | ERROR_vsync
              | ERROR_red | ERROR_green | ERROR_blue | ERROR_x | ERROR_y | ERROR_bmem_addr | ERROR_bmem_color;


    initial begin
        $monitor("#%02d {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h%h, 32'h%h, 32'h%h, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 16'h%h, 1'b%b, 5'b%b, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 5'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 2'b%b, 2'b%b, 1'b%b, 1'b%b, 2'b%b, 1'b%b, 2'b%b};",
                  $time, pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel);
        
        $monitor("#%02d {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h%h, 4'h%h, 1'b%b, 1'b%b, 1'b%b, 1'b%b, 4'h%h, 4'h%h, 4'h%h, 10'h%h, 10'h%h, 12'h%h, 12'h%h};",
                  $time, smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color);

        $monitor("#%02d {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b%b, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h};",
                  $time, sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata);
    end
    
endmodule



// CHECKER MODULE

module selfcheck_nopause();
    logic  [31:0] pc;
    logic  [31:0] instr;
    logic  [31:0] mem_addr;
    logic         mem_wr;
    logic  [31:0] mem_readdata;
    logic  [31:0] mem_writedata;
    logic  [31:0] period;
    logic  [15:0] LED;
    logic         werf;
    logic   [4:0] alufn;
    logic         Z;
    logic  [31:0] ReadData1;
    logic  [31:0] ReadData2;
    logic  [31:0] alu_result;
    logic  [4:0]  reg_writeaddr;
    logic  [31:0] reg_writedata;
    logic  [31:0] signImm;
    logic  [31:0] aluA;
    logic  [31:0] aluB;
    logic   [1:0] pcsel;
    logic   [1:0] wasel;
    logic         sgnext;
    logic         bsel;
    logic   [1:0] wdsel;
    logic         wr;
    logic   [1:0] asel;
    logic  [10:0] smem_addr;
    logic   [3:0] charcode;
    logic dmem_wr;
    logic smem_wr;
    logic hsync;
    logic vsync;
    logic   [3:0] red;
    logic   [3:0] green;
    logic   [3:0] blue;
    logic   [9:0] x;
    logic   [9:0] y;
    logic  [11:0] bmem_addr;
    logic  [11:0] bmem_color;
    logic         sound_wr, lights_wr;
    logic  [31:0] smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata;
    
initial begin
fork

#00 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400000, 32'h3c1d1001, 32'h10010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10010000, 5'h1d, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#00 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h000, 10'h000, 12'h000, 12'hf00};
#00 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'hxxxxxxxx};
#01 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400004, 32'h37bd1000, 32'h10011000, 1'b0, 32'h00000000, 32'h10010000, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'h10010000, 32'h10011000, 5'h1d, 32'h10011000, 32'h00001000, 32'h10010000, 32'h00001000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#01 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000000, 32'h10010000};
#02 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400008, 32'h3c08ffff, 32'hffff0000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'hffff0000, 5'h08, 32'hffff0000, 32'hxxxxffff, 32'h00000010, 32'hxxxxffff, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#02 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hffff0000, 32'h00000000, 32'hxxxxxxxx};
#03 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040000c, 32'h3508ffff, 32'hffffffff, 1'b0, 32'h00000000, 32'hffff0000, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'hffff0000, 32'hffff0000, 32'hffffffff, 5'h08, 32'hffffffff, 32'h0000ffff, 32'hffff0000, 32'h0000ffff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#03 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hffffffff, 32'h00000000, 32'hffff0000};
#04 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400010, 32'h2009ffff, 32'hffffffff, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'hffffffff, 5'h09, 32'hffffffff, 32'hffffffff, 32'h00000000, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#04 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hffffffff, 32'h00000000, 32'hxxxxxxxx};
#04 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h001, 10'h000, 12'h001, 12'hf00};
#05 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h1509003a, 32'h00000000, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h0000003a, 32'hffffffff, 32'hffffffff, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#05 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hffffffff};
#06 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00084600, 32'hff000000, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hffffffff, 32'hff000000, 5'h08, 32'hff000000, 32'h00004600, 32'h00000018, 32'hffffffff, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#06 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff000000, 32'h00000000, 32'hffffffff};
#07 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h3508f000, 32'hff00f000, 1'b0, 32'h00000000, 32'hff000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'hff000000, 32'hff000000, 32'hff00f000, 5'h08, 32'hff00f000, 32'h0000f000, 32'hff000000, 32'h0000f000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#07 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff00f000, 32'h00000000, 32'hff000000};
#08 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h00084203, 32'hffff00f0, 1'b0, 32'h00000000, 32'hff00f000, 32'h00000000, 16'h0000, 1'b1, 5'bx1110, 1'b0, 32'h00000000, 32'hff00f000, 32'hffff00f0, 5'h08, 32'hffff00f0, 32'h00004203, 32'h00000008, 32'hff00f000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#08 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hffff00f0, 32'h00000000, 32'hff00f000};
#08 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h002, 10'h000, 12'h002, 12'hf00};
#09 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h00084102, 32'h0ffff00f, 1'b0, 32'h00000000, 32'hffff00f0, 32'h00000000, 16'h0000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'hffff00f0, 32'h0ffff00f, 5'h08, 32'h0ffff00f, 32'h00004102, 32'h00000004, 32'hffff00f0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#09 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0ffff00f, 32'h00000000, 32'hffff00f0};
#10 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h340a0003, 32'h00000003, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000003, 5'h0a, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#10 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'hxxxxxxxx};
#11 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h01495022, 32'h00000004, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 16'h0000, 1'b1, 5'b1xx01, 1'b0, 32'h00000003, 32'hffffffff, 32'h00000004, 5'h0a, 32'h00000004, 32'h00005022, 32'h00000003, 32'hffffffff, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#11 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000004, 32'h00000000, 32'hffffffff};
#12 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h01484004, 32'hffff00f0, 1'b0, 32'h00000000, 32'h0ffff00f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000004, 32'h0ffff00f, 32'hffff00f0, 5'h08, 32'hffff00f0, 32'h00004004, 32'h00000004, 32'h0ffff00f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#12 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hffff00f0, 32'h00000000, 32'h0ffff00f};
#12 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h003, 10'h000, 12'h003, 12'hf00};
#13 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h01484007, 32'hfffff00f, 1'b0, 32'h00000000, 32'hffff00f0, 32'h00000000, 16'h0000, 1'b1, 5'bx1110, 1'b0, 32'h00000004, 32'hffff00f0, 32'hfffff00f, 5'h08, 32'hfffff00f, 32'h00004007, 32'h00000004, 32'hffff00f0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#13 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hfffff00f, 32'h00000000, 32'hffff00f0};
#14 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h01484006, 32'h0fffff00, 1'b0, 32'h00000000, 32'hfffff00f, 32'h00000000, 16'h0000, 1'b1, 5'bx1010, 1'b0, 32'h00000004, 32'hfffff00f, 32'h0fffff00, 5'h08, 32'h0fffff00, 32'h00004006, 32'h00000004, 32'hfffff00f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#14 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0fffff00, 32'h00000000, 32'hfffff00f};
#15 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h01484004, 32'hfffff000, 1'b0, 32'h00000000, 32'h0fffff00, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000004, 32'h0fffff00, 32'hfffff000, 5'h08, 32'hfffff000, 32'h00004004, 32'h00000004, 32'h0fffff00, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#15 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000000, 32'h00000000, 32'hfffff000, 32'h00000000, 32'h0fffff00};
#16 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h010a582a, 32'h00000001, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'hfffff000, 32'h00000004, 32'h00000001, 5'h0b, 32'h00000001, 32'h0000582a, 32'hfffff000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#16 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000004};
#16 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h004, 10'h000, 12'h004, 12'hf00};
#17 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h010a582b, 32'h00000000, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b1x111, 1'b1, 32'hfffff000, 32'h00000004, 32'h00000000, 5'h0b, 32'h00000000, 32'h0000582b, 32'hfffff000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#17 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000004};
#18 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h20080005, 32'h00000005, 1'b0, 32'h00000000, 32'hfffff000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hfffff000, 32'h00000005, 5'h08, 32'h00000005, 32'h00000005, 32'h00000000, 32'h00000005, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#18 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000005, 32'h00000000, 32'hfffff000};
#19 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h290b000a, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000005, 32'h00000000, 32'h00000001, 5'h0b, 32'h00000001, 32'h0000000a, 32'h00000005, 32'h0000000a, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#19 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#20 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h2d0b0004, 32'h00000000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x111, 1'b1, 32'h00000005, 32'h00000001, 32'h00000000, 5'h0b, 32'h00000000, 32'h00000004, 32'h00000005, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#20 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001};
#20 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h005, 10'h000, 12'h005, 12'hf00};
#21 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h2008fffb, 32'hfffffffb, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000005, 32'hfffffffb, 5'h08, 32'hfffffffb, 32'hfffffffb, 32'h00000000, 32'hfffffffb, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#21 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hfffffffb, 32'h00000000, 32'h00000005};
#22 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h2d0b0005, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b1x111, 1'b1, 32'hfffffffb, 32'h00000000, 32'h00000000, 5'h0b, 32'h00000000, 32'h00000005, 32'hfffffffb, 32'h00000005, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#22 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#23 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h20080014, 32'h00000014, 1'b0, 32'h00000000, 32'hfffffffb, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hfffffffb, 32'h00000014, 5'h08, 32'h00000014, 32'h00000014, 32'h00000000, 32'h00000014, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#23 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000014, 32'h00000000, 32'hfffffffb};
#24 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400060, 32'h2d0bffff, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b1x111, 1'b0, 32'h00000014, 32'h00000000, 32'h00000001, 5'h0b, 32'h00000001, 32'hffffffff, 32'h00000014, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#24 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#24 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h006, 10'h000, 12'h006, 12'hf00};
#25 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400064, 32'h3c0b1010, 32'h10100000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10100000, 5'h0b, 32'h10100000, 32'h00001010, 32'h00000010, 32'h00001010, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#25 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10100000, 32'h00000000, 32'h00000001};
#26 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400068, 32'h356b1010, 32'h10101010, 1'b0, 32'h00000000, 32'h10100000, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10100000, 32'h10100000, 32'h10101010, 5'h0b, 32'h10101010, 32'h00001010, 32'h10100000, 32'h00001010, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#26 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10101010, 32'h00000000, 32'h10100000};
#27 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040006c, 32'h3c0c0101, 32'h01010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h01010000, 5'h0c, 32'h01010000, 32'h00000101, 32'h00000010, 32'h00000101, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#27 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h01010000, 32'h00000000, 32'hxxxxxxxx};
#28 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400070, 32'h218c1010, 32'h01011010, 1'b0, 32'hxxxxxxxx, 32'h01010000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h01010000, 32'h01010000, 32'h01011010, 5'h0c, 32'h01011010, 32'h00001010, 32'h01010000, 32'h00001010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#28 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h01011010, 32'hxxxxxxxx, 32'h01010000};
#28 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h007, 10'h000, 12'h007, 12'hf00};
#29 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h318dffff, 32'h00001010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0000, 1'b0, 32'h01011010, 32'hxxxxxxxx, 32'h00001010, 5'h0d, 32'h00001010, 32'h0000ffff, 32'h01011010, 32'h0000ffff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#29 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00001010, 32'h00000000, 32'hxxxxxxxx};
#30 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h39adffff, 32'h0000efef, 1'b0, 32'h00000000, 32'h00001010, 32'h00000000, 16'h0000, 1'b1, 5'bx1000, 1'b0, 32'h00001010, 32'h00001010, 32'h0000efef, 5'h0d, 32'h0000efef, 32'h0000ffff, 32'h00001010, 32'h0000ffff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#30 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000efef, 32'h00000000, 32'h00001010};
#31 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040007c, 32'h016c6824, 32'h00001010, 1'b0, 32'h00000000, 32'h01011010, 32'h00000000, 16'h0000, 1'b1, 5'bx0000, 1'b0, 32'h10101010, 32'h01011010, 32'h00001010, 5'h0d, 32'h00001010, 32'h00006824, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#31 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00001010, 32'h00000000, 32'h01011010};
#32 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400080, 32'h016c6825, 32'h11111010, 1'b0, 32'hxxxxxxxx, 32'h01011010, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10101010, 32'h01011010, 32'h11111010, 5'h0d, 32'h11111010, 32'h00006825, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#32 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h008, 10'h000, 12'h008, 12'hf00};
#32 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h11111010, 32'hxxxxxxxx, 32'h01011010};
#33 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400084, 32'h016c6826, 32'h11110000, 1'b0, 32'h00000000, 32'h01011010, 32'h00000000, 16'h0000, 1'b1, 5'bx1000, 1'b0, 32'h10101010, 32'h01011010, 32'h11110000, 5'h0d, 32'h11110000, 32'h00006826, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#33 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h11110000, 32'h00000000, 32'h01011010};
#34 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400088, 32'h016c6827, 32'heeeeefef, 1'b0, 32'h00000003, 32'h01011010, 32'h00000000, 16'h0000, 1'b1, 5'bx1100, 1'b0, 32'h10101010, 32'h01011010, 32'heeeeefef, 5'h0d, 32'heeeeefef, 32'h00006827, 32'h10101010, 32'h01011010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#34 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'heeeeefef, 32'h00000003, 32'h01011010};
#35 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040008c, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#35 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'hxxxxxxxx};
#36 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'h00200821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#36 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'h00000000};
#36 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h009, 10'h000, 12'h009, 12'hf00};
#37 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h8c240004, 32'h10010004, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010004, 5'h04, 32'h00000003, 32'h00000004, 32'h10010000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#37 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h10010004, 32'h00000003, 32'hxxxxxxxx};
#38 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400098, 32'h20840002, 32'h00000005, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000005, 5'h04, 32'h00000005, 32'h00000002, 32'h00000003, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#38 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000005, 32'h00000000, 32'h00000003};
#39 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040009c, 32'h2484fffe, 32'h00000003, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000003, 5'h04, 32'h00000003, 32'hfffffffe, 32'h00000005, 32'hfffffffe, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#39 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000005};
#40 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000a0, 32'h3c010040, 32'h00400000, 1'b0, 32'h00000000, 32'h10010000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h00400000, 5'h01, 32'h00400000, 32'h00000040, 32'h00000010, 32'h00000040, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#40 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00400000, 32'h00000000, 32'h10010000};
#40 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00a, 10'h000, 12'h00a, 12'hf00};
#41 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000a4, 32'h34300104, 32'h00400104, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h00400000, 32'hxxxxxxxx, 32'h00400104, 5'h10, 32'h00400104, 32'h00000104, 32'h00400000, 32'h00000104, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#41 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00400104, 32'h00000000, 32'hxxxxxxxx};
#42 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000a8, 32'h0200f809, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00400104, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h004000ac, 32'hxxxxf809, 32'hxxxxxxxx, 32'hxxxxxX0X, 2'b11, 2'b00, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#42 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#43 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'h23bdfff8, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff8, 5'h1d, 32'h10010ff8, 32'hfffffff8, 32'h10011000, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#43 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'hxxxxxxxx, 32'h10011000};
#44 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafbf0004, 32'h10010ffc, 1'b1, 32'hxxxxxxxx, 32'h004000ac, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h004000ac, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff8, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#44 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'hxxxxxxxx, 32'h004000ac};
#44 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00b, 10'h000, 12'h00b, 12'hf00};
#45 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'hxxxxxxxx, 32'h00000003};
#45 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'hafa40000, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h00000003, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#46 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000014};
#46 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h28880002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000014, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b1, 32'h00000003, 32'h00000014, 32'h00000000, 5'h08, 32'h00000000, 32'h00000002, 32'h00000003, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#46 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00b, 10'h000, 12'h00b, 12'hf00};
#47 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h11000002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#47 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#48 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h2084ffff, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'hffffffff, 32'h00000003, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#48 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h000, 12'h00c, 12'hf00};
#48 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#49 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h0c100041, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h00400128, 32'h00000041, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#49 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#50 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'h23bdfff8, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10010ff8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h10010ff8, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff8, 32'h10010ff8, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#50 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8};
#51 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafbf0004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'h00400128, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400128, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#51 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hxxxxxxxx, 32'h00400128};
#51 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00c, 10'h000, 12'h00c, 12'hf00};
#52 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000002};
#52 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'hafa40000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000002, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#52 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00d, 10'h000, 12'h00d, 12'hf00};
#53 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#53 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h28880002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b1, 32'h00000002, 32'h00000000, 32'h00000000, 5'h08, 32'h00000000, 32'h00000002, 32'h00000002, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#53 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00d, 10'h000, 12'h00d, 12'hf00};
#54 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h11000002, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#55 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h2084ffff, 32'h00000001, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000002, 32'h00000002, 32'h00000001, 5'h04, 32'h00000001, 32'hffffffff, 32'h00000002, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#55 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000002};
#56 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h0c100041, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h00400128, 32'h00000041, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#56 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#56 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00e, 10'h000, 12'h00e, 12'hf00};
#57 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'h23bdfff8, 32'h10010fe8, 1'b0, 32'hxxxxxxxx, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10010fe8, 5'h1d, 32'h10010fe8, 32'hfffffff8, 32'h10010ff0, 32'hfffffff8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#57 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010fe8, 32'hxxxxxxxx, 32'h10010ff0};
#58 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafbf0004, 32'h10010fec, 1'b1, 32'hxxxxxxxx, 32'h00400128, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010fe8, 32'h00400128, 32'h10010fec, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010fe8, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#58 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010fec, 32'hxxxxxxxx, 32'h00400128};
#58 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00e, 10'h000, 12'h00e, 12'hf00};
#59 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10010fe8, 32'hxxxxxxxx, 32'h00000001};
#59 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'hafa40000, 32'h10010fe8, 1'b1, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010fe8, 32'h00000001, 32'h10010fe8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010fe8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#60 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#60 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h28880002, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'h08, 32'h00000001, 32'h00000002, 32'h00000001, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#60 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h000, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h00f, 10'h000, 12'h00f, 12'hf00};
#61 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h11000002, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'h00000002, 32'h00000001, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#62 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h00041020, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000001, 5'h02, 32'h00000001, 32'h00001020, 32'h00000000, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#62 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#63 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h0810004e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h0000004e, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#63 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#64 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fbf0004, 32'h10010fec, 1'b0, 32'h00400128, 32'h00400128, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010fe8, 32'h00400128, 32'h10010fec, 5'h1f, 32'h00400128, 32'h00000004, 32'h10010fe8, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#64 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h010, 10'h000, 12'h000, 12'hf00};
#64 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00400128, 32'h00000000, 32'h00000000, 32'h10010fec, 32'h00400128, 32'h00400128};
#65 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h23bd0008, 32'h10010ff0, 1'b0, 32'h00000002, 32'h10010fe8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010fe8, 32'h10010fe8, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'h00000008, 32'h10010fe8, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#65 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000002, 32'h10010fe8};
#66 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400128, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#66 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#67 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h8fa40000, 32'h10010ff0, 1'b0, 32'h00000002, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff0, 5'h04, 32'h00000002, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#67 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000002, 32'h00000001};
#68 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'h00441020, 32'h00000003, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000002, 32'h00000003, 5'h02, 32'h00000003, 32'h00001020, 32'h00000001, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#68 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000002};
#68 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h011, 10'h000, 12'h001, 12'hf00};
#69 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h00441020, 32'h00000005, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000002, 32'h00000005, 5'h02, 32'h00000005, 32'h00001020, 32'h00000003, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#69 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000005, 32'h00000000, 32'h00000002};
#70 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h2042ffff, 32'h00000004, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000004, 5'h02, 32'h00000004, 32'hffffffff, 32'h00000005, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#70 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000005};
#71 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fbf0004, 32'h10010ff4, 1'b0, 32'h00400128, 32'h00400128, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400128, 32'h10010ff4, 5'h1f, 32'h00400128, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#71 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400128, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'h00400128, 32'h00400128};
#72 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h23bd0008, 32'h10010ff8, 1'b0, 32'h00000003, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10010ff8, 5'h1d, 32'h10010ff8, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#72 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h012, 10'h000, 12'h002, 12'hf00};
#72 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000003, 32'h10010ff0};
#73 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400128, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#73 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#74 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h8fa40000, 32'h10010ff8, 1'b0, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h00000002, 32'h10010ff8, 5'h04, 32'h00000003, 32'h00000000, 32'h10010ff8, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#74 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000003, 32'h00000002};
#75 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'h00441020, 32'h00000007, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000003, 32'h00000007, 5'h02, 32'h00000007, 32'h00001020, 32'h00000004, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#75 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000007, 32'h00000000, 32'h00000003};
#76 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h00441020, 32'h0000000a, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000007, 32'h00000003, 32'h0000000a, 5'h02, 32'h0000000a, 32'h00001020, 32'h00000007, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#76 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000a, 32'h00000000, 32'h00000003};
#76 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h013, 10'h000, 12'h003, 12'hf00};
#77 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h2042ffff, 32'h00000009, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000a, 32'h0000000a, 32'h00000009, 5'h02, 32'h00000009, 32'hffffffff, 32'h0000000a, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#77 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000009, 32'h00000000, 32'h0000000a};
#78 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fbf0004, 32'h10010ffc, 1'b0, 32'h004000ac, 32'h00400128, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h00400128, 32'h10010ffc, 5'h1f, 32'h004000ac, 32'h00000004, 32'h10010ff8, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#78 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000ac, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000ac, 32'h00400128};
#79 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h23bd0008, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff8, 32'h10010ff8, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000008, 32'h10010ff8, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#79 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000000, 32'h10010ff8};
#80 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000ac, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#80 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#80 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h014, 10'h000, 12'h004, 12'hf00};
#81 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ac, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00400000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00400000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#81 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'h00400000};
#82 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b0, 32'h00200821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#82 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'h00000000};
#83 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b4, 32'hac220000, 32'h10010000, 1'b1, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000009, 32'h10010000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#83 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'h00000009};
#83 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h014, 10'h000, 12'h004, 12'hf00};
#84 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000003e8, 32'h00000000, 32'h00000003};
#84 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b8, 32'h200403e8, 32'h000003e8, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h000003e8, 5'h04, 32'h000003e8, 32'h000003e8, 32'h00000000, 32'h000003e8, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#84 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h015, 10'h000, 12'h005, 12'hf00};
#85 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000bc, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#85 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#86 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c0, 32'h24050000, 32'h00000000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 5'h05, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#86 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hxxxxxxxx};
#87 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c4, 32'h24060000, 32'h00000000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 5'h06, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#88 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h000003e8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h000003e8, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#88 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h000003e8};
#88 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h016, 10'h000, 12'h006, 12'hf00};
#89 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#89 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#90 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000002, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#90 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000002, 32'h10011000};
#91 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000ac, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#91 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000ac, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000ac, 32'h004000d0};
#91 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h016, 10'h000, 12'h006, 12'hf00};
#92 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000003, 32'h00000001};
#92 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#92 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h017, 10'h000, 12'h007, 12'hf00};
#93 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400128, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'h00400128, 32'hffffffff};
#93 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'h00400128, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#94 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000002, 32'h00000004};
#94 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000002, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#95 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000000, 32'h10010000};
#95 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h10010000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#95 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h017, 10'h000, 12'h007, 12'hf00};
#96 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#96 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000000, 32'h00000001};
#96 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h018, 10'h000, 12'h008, 12'hf00};
#97 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004940, 32'h00000005, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#97 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#98 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h0a, 32'h00000000, 32'h000050c0, 32'h00000003, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#99 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#100 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#100 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h019, 10'h000, 12'h009, 12'hf00};
#101 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004880, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#102 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000000, 32'h10020000, 5'h08, 32'h10020000, 32'h00004020, 32'h10020000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#102 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000000, 32'h00000000};
#103 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020000, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000002, 32'h10020000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#103 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000000, 32'h00000002};
#103 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h019, 10'h000, 12'h009, 12'hf00};
#104 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#104 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#104 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01a, 10'h000, 12'h00a, 12'hf00};
#105 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020000, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#105 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020000};
#106 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000000, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#106 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000000};
#107 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000000, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#107 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000000};
#108 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#108 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#108 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01b, 10'h000, 12'h00b, 12'hf00};
#109 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#109 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#110 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#110 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#111 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#111 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#112 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#112 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01c, 10'h000, 12'h00c, 12'hf00};
#112 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#113 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#113 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#114 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#114 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#115 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#115 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#115 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01c, 10'h000, 12'h00c, 12'hf00};
#116 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#116 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#116 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01d, 10'h000, 12'h00d, 12'hf00};
#117 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#117 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#118 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#118 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#119 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000002, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#119 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000002, 32'h10020000};
#119 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01d, 10'h000, 12'h00d, 12'hf00};
#120 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000002, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#120 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01e, 10'h000, 12'h00e, 12'hf00};
#120 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000002, 32'h00000001};
#121 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004940, 32'h00000005, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#121 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#122 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h0a, 32'h00000000, 32'h000050c0, 32'h00000003, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#123 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#124 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004820, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#124 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01f, 10'h000, 12'h00f, 12'hf00};
#125 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h09, 32'h00000000, 32'h00004880, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#126 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020000, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000000, 32'h10020000, 5'h08, 32'h10020000, 32'h00004020, 32'h10020000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#126 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000002, 32'h00000000};
#127 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020000, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000003, 32'h10020000, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#127 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000002, 32'h00000003};
#127 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h001, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h01f, 10'h000, 12'h00f, 12'hf00};
#128 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#128 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#128 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h020, 10'h000, 12'h000, 12'hf00};
#129 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020000, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#129 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020000};
#130 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000000, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#130 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000000};
#131 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000000, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#131 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000000};
#132 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#132 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#132 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h021, 10'h000, 12'h001, 12'hf00};
#133 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#133 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#134 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000001, 5'h05, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#134 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#135 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000001, 5'h06, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#136 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000001, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000001, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#136 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#136 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h022, 10'h000, 12'h002, 12'hf00};
#137 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#137 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#138 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#138 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#139 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#139 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#140 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#140 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h023, 10'h000, 12'h003, 12'hf00};
#140 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#141 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#141 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#141 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h023, 10'h000, 12'h003, 12'hf00};
#142 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#142 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#143 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#143 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#144 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#144 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h000, 12'h004, 12'hf00};
#144 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#145 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#145 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#145 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h024, 10'h000, 12'h004, 12'hf00};
#146 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#146 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#147 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000020, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000020, 5'h09, 32'h00000020, 32'h00004940, 32'h00000005, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#147 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000020, 32'h00000000, 32'h00000001};
#148 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000008, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000008, 5'h0a, 32'h00000008, 32'h000050c0, 32'h00000003, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#148 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h025, 10'h000, 12'h005, 12'hf00};
#148 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000008, 32'h00000000, 32'h00000001};
#149 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000028, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000020, 32'h00000008, 32'h00000028, 5'h09, 32'h00000028, 32'h00004820, 32'h00000020, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#149 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000028, 32'h00000000, 32'h00000008};
#150 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000029, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000028, 32'h00000001, 32'h00000029, 5'h09, 32'h00000029, 32'h00004820, 32'h00000028, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#150 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000029, 32'h00000000, 32'h00000001};
#151 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000029, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000029, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004880, 32'h00000002, 32'h00000029, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#151 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a4, 32'h00000000, 32'h00000029};
#152 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100200a4, 1'b0, 32'h00000001, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000000a4, 32'h100200a4, 5'h08, 32'h100200a4, 32'h00004020, 32'h10020000, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#152 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100200a4, 32'h00000001, 32'h000000a4};
#152 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h000, 12'h006, 12'hf00};
#153 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100200a4, 1'b1, 32'h00000001, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100200a4, 32'h00000002, 32'h100200a4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100200a4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#153 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100200a4, 32'h00000001, 32'h00000002};
#153 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h000, 12'h006, 12'hf00};
#154 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#154 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#154 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h026, 10'h000, 12'h006, 12'hf00};
#155 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100200a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100200a4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#155 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100200a4};
#156 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000000a4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#156 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000000a4};
#156 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h027, 10'h000, 12'h007, 12'hf00};
#157 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000008, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#157 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000008};
#158 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#158 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#159 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#159 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#160 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#160 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h028, 10'h000, 12'h008, 12'hf00};
#160 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#161 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#161 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#162 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#162 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#163 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#163 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#164 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#164 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h029, 10'h000, 12'h009, 12'hf00};
#164 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#165 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#165 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#165 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h029, 10'h000, 12'h009, 12'hf00};
#166 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#166 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#167 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#167 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#168 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#168 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02a, 10'h000, 12'h00a, 12'hf00};
#168 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#169 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#169 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#169 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02a, 10'h000, 12'h00a, 12'hf00};
#170 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#170 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#171 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000020, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000020, 5'h09, 32'h00000020, 32'h00004940, 32'h00000005, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#171 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000020, 32'h00000000, 32'h00000001};
#172 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000008, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000008, 5'h0a, 32'h00000008, 32'h000050c0, 32'h00000003, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#172 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02b, 10'h000, 12'h00b, 12'hf00};
#172 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000008, 32'h00000000, 32'h00000001};
#173 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000028, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000020, 32'h00000008, 32'h00000028, 5'h09, 32'h00000028, 32'h00004820, 32'h00000020, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#173 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000028, 32'h00000000, 32'h00000008};
#174 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000029, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000028, 32'h00000001, 32'h00000029, 5'h09, 32'h00000029, 32'h00004820, 32'h00000028, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#174 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000029, 32'h00000000, 32'h00000001};
#175 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000029, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000029, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004880, 32'h00000002, 32'h00000029, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#175 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a4, 32'h00000000, 32'h00000029};
#176 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100200a4, 1'b0, 32'h00000002, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000000a4, 32'h100200a4, 5'h08, 32'h100200a4, 32'h00004020, 32'h10020000, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#176 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100200a4, 32'h00000002, 32'h000000a4};
#176 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h000, 12'h00c, 12'hf00};
#177 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100200a4, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100200a4, 32'h00000003, 32'h100200a4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100200a4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#177 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100200a4, 32'h00000002, 32'h00000003};
#177 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h000, 12'h00c, 12'hf00};
#178 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#178 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#178 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02c, 10'h000, 12'h00c, 12'hf00};
#179 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100200a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100200a4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#179 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100200a4};
#180 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000000a4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#180 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000000a4};
#180 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02d, 10'h000, 12'h00d, 12'hf00};
#181 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000008, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#181 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000008};
#182 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#182 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#183 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#183 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#184 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000002, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000001, 32'h00000002, 5'h05, 32'h00000002, 32'h00000001, 32'h00000001, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#184 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02e, 10'h000, 12'h00e, 12'hf00};
#184 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000001};
#185 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000002, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000001, 32'h00000001, 32'h00000002, 5'h06, 32'h00000002, 32'h00000001, 32'h00000001, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#186 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000002, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000002, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#186 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#187 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#187 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#188 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#188 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02f, 10'h000, 12'h00f, 12'hf00};
#188 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#189 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#189 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#190 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#190 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#191 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#191 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#191 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h002, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h02f, 10'h000, 12'h00f, 12'hf00};
#192 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#192 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#192 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h030, 10'h000, 12'h100, 12'h0f0};
#193 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#193 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#194 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#194 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#195 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#195 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#195 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h030, 10'h000, 12'h100, 12'h0f0};
#196 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#196 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h031, 10'h000, 12'h101, 12'h0f0};
#196 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#197 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000040, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000040, 5'h09, 32'h00000040, 32'h00004940, 32'h00000005, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#197 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000040, 32'h00000000, 32'h00000002};
#198 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000010, 5'h0a, 32'h00000010, 32'h000050c0, 32'h00000003, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#198 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000010, 32'h00000000, 32'h00000002};
#199 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000050, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000040, 32'h00000010, 32'h00000050, 5'h09, 32'h00000050, 32'h00004820, 32'h00000040, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#199 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000050, 32'h00000000, 32'h00000010};
#200 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000052, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000050, 32'h00000002, 32'h00000052, 5'h09, 32'h00000052, 32'h00004820, 32'h00000050, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#200 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000052, 32'h00000000, 32'h00000002};
#200 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h032, 10'h000, 12'h102, 12'h0f0};
#201 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000148, 1'b0, 32'h00000000, 32'h00000052, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000052, 32'h00000148, 5'h09, 32'h00000148, 32'h00004880, 32'h00000002, 32'h00000052, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#201 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000148, 32'h00000000, 32'h00000052};
#202 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020148, 1'b0, 32'h00000003, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000148, 32'h10020148, 5'h08, 32'h10020148, 32'h00004020, 32'h10020000, 32'h00000148, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#202 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020148, 32'h00000003, 32'h00000148};
#203 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020148, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020148, 32'h00000002, 32'h10020148, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020148, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#203 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020148, 32'h00000003, 32'h00000002};
#203 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h032, 10'h000, 12'h102, 12'h0f0};
#204 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#204 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#204 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h033, 10'h000, 12'h103, 12'h0f0};
#205 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020148, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#205 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020148};
#206 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000148, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#206 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000148};
#207 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#207 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000010};
#208 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#208 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#208 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h034, 10'h000, 12'h104, 12'h0f0};
#209 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#209 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#210 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#210 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#211 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#211 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#212 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#212 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h035, 10'h000, 12'h105, 12'h0f0};
#212 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#213 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#213 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#214 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#214 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#215 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#215 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#215 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h035, 10'h000, 12'h105, 12'h0f0};
#216 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#216 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#216 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h036, 10'h000, 12'h106, 12'h0f0};
#217 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#217 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#218 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#218 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#219 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#219 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#219 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h036, 10'h000, 12'h106, 12'h0f0};
#220 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#220 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h037, 10'h000, 12'h107, 12'h0f0};
#220 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#221 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000040, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000040, 5'h09, 32'h00000040, 32'h00004940, 32'h00000005, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#221 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000040, 32'h00000000, 32'h00000002};
#222 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000002, 32'h00000010, 5'h0a, 32'h00000010, 32'h000050c0, 32'h00000003, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#222 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000010, 32'h00000000, 32'h00000002};
#223 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000050, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000040, 32'h00000010, 32'h00000050, 5'h09, 32'h00000050, 32'h00004820, 32'h00000040, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#223 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000050, 32'h00000000, 32'h00000010};
#224 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000052, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000050, 32'h00000002, 32'h00000052, 5'h09, 32'h00000052, 32'h00004820, 32'h00000050, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#224 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000052, 32'h00000000, 32'h00000002};
#224 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h038, 10'h000, 12'h108, 12'h0f0};
#225 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000148, 1'b0, 32'h00000000, 32'h00000052, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000052, 32'h00000148, 5'h09, 32'h00000148, 32'h00004880, 32'h00000002, 32'h00000052, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#225 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000148, 32'h00000000, 32'h00000052};
#226 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020148, 1'b0, 32'h00000002, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000148, 32'h10020148, 5'h08, 32'h10020148, 32'h00004020, 32'h10020000, 32'h00000148, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#226 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020148, 32'h00000002, 32'h00000148};
#227 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020148, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020148, 32'h00000003, 32'h10020148, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020148, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#227 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020148, 32'h00000002, 32'h00000003};
#227 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h038, 10'h000, 12'h108, 12'h0f0};
#228 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#228 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#228 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h039, 10'h000, 12'h109, 12'h0f0};
#229 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020148, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#229 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020148};
#230 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000148, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#230 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000148};
#231 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#231 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000010};
#232 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#232 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#232 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03a, 10'h000, 12'h10a, 12'h0f0};
#233 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#233 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#234 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000003, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000002, 32'h00000002, 32'h00000003, 5'h05, 32'h00000003, 32'h00000001, 32'h00000002, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#234 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000002};
#235 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000003, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000002, 32'h00000002, 32'h00000003, 5'h06, 32'h00000003, 32'h00000001, 32'h00000002, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#236 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000003, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000003, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#236 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#236 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03b, 10'h000, 12'h10b, 12'h0f0};
#237 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#237 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#238 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#238 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#239 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#239 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#240 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#240 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03c, 10'h000, 12'h10c, 12'h0f0};
#240 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#241 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#241 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#241 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03c, 10'h000, 12'h10c, 12'h0f0};
#242 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#242 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#243 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#243 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#244 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#244 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03d, 10'h000, 12'h10d, 12'h0f0};
#244 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#245 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#245 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#245 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03d, 10'h000, 12'h10d, 12'h0f0};
#246 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#246 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#247 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000060, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000003, 32'h00000060, 5'h09, 32'h00000060, 32'h00004940, 32'h00000005, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#247 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000060, 32'h00000000, 32'h00000003};
#248 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000018, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000003, 32'h00000018, 5'h0a, 32'h00000018, 32'h000050c0, 32'h00000003, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#248 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03e, 10'h000, 12'h10e, 12'h0f0};
#248 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000018, 32'h00000000, 32'h00000003};
#249 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000078, 1'b0, 32'h00000000, 32'h00000018, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000060, 32'h00000018, 32'h00000078, 5'h09, 32'h00000078, 32'h00004820, 32'h00000060, 32'h00000018, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#249 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000078, 32'h00000000, 32'h00000018};
#250 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000007b, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000078, 32'h00000003, 32'h0000007b, 5'h09, 32'h0000007b, 32'h00004820, 32'h00000078, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#250 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000007b, 32'h00000000, 32'h00000003};
#251 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000001ec, 1'b0, 32'h00000000, 32'h0000007b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000007b, 32'h000001ec, 5'h09, 32'h000001ec, 32'h00004880, 32'h00000002, 32'h0000007b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#251 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001ec, 32'h00000000, 32'h0000007b};
#252 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100201ec, 1'b0, 32'h00000001, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000001ec, 32'h100201ec, 5'h08, 32'h100201ec, 32'h00004020, 32'h10020000, 32'h000001ec, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#252 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100201ec, 32'h00000001, 32'h000001ec};
#252 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03f, 10'h000, 12'h10f, 12'h0f0};
#253 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100201ec, 1'b1, 32'h00000001, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100201ec, 32'h00000002, 32'h100201ec, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100201ec, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#253 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100201ec, 32'h00000001, 32'h00000002};
#253 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03f, 10'h000, 12'h10f, 12'h0f0};
#254 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#254 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#254 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h003, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h03f, 10'h000, 12'h10f, 12'h0f0};
#255 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100201ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100201ec, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#255 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100201ec};
#256 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000001ec, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#256 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000001ec};
#256 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h040, 10'h000, 12'h100, 12'h0f0};
#257 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000018, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000018, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#257 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000018};
#258 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#258 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#259 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#259 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#260 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#260 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h041, 10'h000, 12'h101, 12'h0f0};
#260 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#261 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#261 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#262 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#262 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#263 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#263 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#264 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#264 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h042, 10'h000, 12'h102, 12'h0f0};
#264 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#265 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#265 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#265 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h042, 10'h000, 12'h102, 12'h0f0};
#266 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#266 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#267 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#267 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#268 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#268 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h043, 10'h000, 12'h103, 12'h0f0};
#268 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#269 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#269 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#269 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h043, 10'h000, 12'h103, 12'h0f0};
#270 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#270 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#271 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000060, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000003, 32'h00000060, 5'h09, 32'h00000060, 32'h00004940, 32'h00000005, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#271 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000060, 32'h00000000, 32'h00000003};
#272 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000018, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000003, 32'h00000018, 5'h0a, 32'h00000018, 32'h000050c0, 32'h00000003, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#272 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h044, 10'h000, 12'h104, 12'h0f0};
#272 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000018, 32'h00000000, 32'h00000003};
#273 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000078, 1'b0, 32'h00000000, 32'h00000018, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000060, 32'h00000018, 32'h00000078, 5'h09, 32'h00000078, 32'h00004820, 32'h00000060, 32'h00000018, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#273 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000078, 32'h00000000, 32'h00000018};
#274 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000007b, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000078, 32'h00000003, 32'h0000007b, 5'h09, 32'h0000007b, 32'h00004820, 32'h00000078, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#274 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000007b, 32'h00000000, 32'h00000003};
#275 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000001ec, 1'b0, 32'h00000000, 32'h0000007b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000007b, 32'h000001ec, 5'h09, 32'h000001ec, 32'h00004880, 32'h00000002, 32'h0000007b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#275 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001ec, 32'h00000000, 32'h0000007b};
#276 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100201ec, 1'b0, 32'h00000002, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000001ec, 32'h100201ec, 5'h08, 32'h100201ec, 32'h00004020, 32'h10020000, 32'h000001ec, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#276 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100201ec, 32'h00000002, 32'h000001ec};
#276 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h045, 10'h000, 12'h105, 12'h0f0};
#277 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100201ec, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100201ec, 32'h00000003, 32'h100201ec, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100201ec, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#277 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100201ec, 32'h00000002, 32'h00000003};
#277 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h045, 10'h000, 12'h105, 12'h0f0};
#278 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#278 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#278 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h045, 10'h000, 12'h105, 12'h0f0};
#279 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100201ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100201ec, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#279 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100201ec};
#280 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000001ec, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#280 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000001ec};
#280 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h046, 10'h000, 12'h106, 12'h0f0};
#281 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000018, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000018, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#281 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000018};
#282 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#282 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#283 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#283 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#284 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000004, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000004, 5'h05, 32'h00000004, 32'h00000001, 32'h00000003, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#284 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h047, 10'h000, 12'h107, 12'h0f0};
#284 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000003};
#285 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000004, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000003, 32'h00000003, 32'h00000004, 5'h06, 32'h00000004, 32'h00000001, 32'h00000003, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#286 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000004, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#286 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#287 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#287 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#288 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#288 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h048, 10'h000, 12'h108, 12'h0f0};
#288 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#289 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#289 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#290 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#290 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#291 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#291 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#291 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h048, 10'h000, 12'h108, 12'h0f0};
#292 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#292 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#292 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h049, 10'h000, 12'h109, 12'h0f0};
#293 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#293 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#294 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#294 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#295 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#295 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#295 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h049, 10'h000, 12'h109, 12'h0f0};
#296 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#296 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04a, 10'h000, 12'h10a, 12'h0f0};
#296 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#297 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000080, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000080, 5'h09, 32'h00000080, 32'h00004940, 32'h00000005, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#297 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000080, 32'h00000000, 32'h00000004};
#298 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000020, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000020, 5'h0a, 32'h00000020, 32'h000050c0, 32'h00000003, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#298 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000020, 32'h00000000, 32'h00000004};
#299 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000a0, 1'b0, 32'h00000000, 32'h00000020, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000080, 32'h00000020, 32'h000000a0, 5'h09, 32'h000000a0, 32'h00004820, 32'h00000080, 32'h00000020, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#299 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a0, 32'h00000000, 32'h00000020};
#300 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000a0, 32'h00000004, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004820, 32'h000000a0, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#300 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a4, 32'h00000000, 32'h00000004};
#300 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04b, 10'h000, 12'h10b, 12'h0f0};
#301 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000290, 1'b0, 32'h00000000, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000a4, 32'h00000290, 5'h09, 32'h00000290, 32'h00004880, 32'h00000002, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#301 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000290, 32'h00000000, 32'h000000a4};
#302 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020290, 1'b0, 32'h00000002, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000290, 32'h10020290, 5'h08, 32'h10020290, 32'h00004020, 32'h10020000, 32'h00000290, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#302 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020290, 32'h00000002, 32'h00000290};
#303 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020290, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020290, 32'h00000002, 32'h10020290, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020290, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#303 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020290, 32'h00000002, 32'h00000002};
#303 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04b, 10'h000, 12'h10b, 12'h0f0};
#304 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#304 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04c, 10'h000, 12'h10c, 12'h0f0};
#304 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#305 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020290, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#305 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020290};
#306 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000290, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#306 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000290};
#307 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000020, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000020, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#307 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000020};
#308 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#308 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#308 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04d, 10'h000, 12'h10d, 12'h0f0};
#309 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#309 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#310 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#310 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#311 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#311 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#312 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#312 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04e, 10'h000, 12'h10e, 12'h0f0};
#312 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#313 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#313 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#314 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#314 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#315 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#315 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#315 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04e, 10'h000, 12'h10e, 12'h0f0};
#316 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#316 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#316 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04f, 10'h000, 12'h10f, 12'h0f0};
#317 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#317 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#318 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#318 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#319 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#319 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#319 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h004, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h04f, 10'h000, 12'h10f, 12'h0f0};
#320 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#320 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h050, 10'h000, 12'h100, 12'h0f0};
#320 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#321 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000080, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000080, 5'h09, 32'h00000080, 32'h00004940, 32'h00000005, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#321 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000080, 32'h00000000, 32'h00000004};
#322 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000020, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000020, 5'h0a, 32'h00000020, 32'h000050c0, 32'h00000003, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#322 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000020, 32'h00000000, 32'h00000004};
#323 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000a0, 1'b0, 32'h00000000, 32'h00000020, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000080, 32'h00000020, 32'h000000a0, 5'h09, 32'h000000a0, 32'h00004820, 32'h00000080, 32'h00000020, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#323 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a0, 32'h00000000, 32'h00000020};
#324 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000a4, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000a0, 32'h00000004, 32'h000000a4, 5'h09, 32'h000000a4, 32'h00004820, 32'h000000a0, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#324 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a4, 32'h00000000, 32'h00000004};
#324 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h051, 10'h000, 12'h101, 12'h0f0};
#325 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000290, 1'b0, 32'h00000000, 32'h000000a4, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000a4, 32'h00000290, 5'h09, 32'h00000290, 32'h00004880, 32'h00000002, 32'h000000a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#325 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000290, 32'h00000000, 32'h000000a4};
#326 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020290, 1'b0, 32'h00000002, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000290, 32'h10020290, 5'h08, 32'h10020290, 32'h00004020, 32'h10020000, 32'h00000290, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#326 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020290, 32'h00000002, 32'h00000290};
#327 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020290, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020290, 32'h00000003, 32'h10020290, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020290, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#327 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020290, 32'h00000002, 32'h00000003};
#327 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h051, 10'h000, 12'h101, 12'h0f0};
#328 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#328 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#328 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h052, 10'h000, 12'h102, 12'h0f0};
#329 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020290, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#329 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020290};
#330 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000290, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#330 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000290};
#331 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000020, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000020, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#331 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000020};
#332 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#332 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#332 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h053, 10'h000, 12'h103, 12'h0f0};
#333 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#333 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#334 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000005, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000005, 5'h05, 32'h00000005, 32'h00000001, 32'h00000004, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#334 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000005, 32'h00000000, 32'h00000004};
#335 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000005, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000005, 5'h06, 32'h00000005, 32'h00000001, 32'h00000004, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#336 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000005, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000005, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#336 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#336 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h054, 10'h000, 12'h104, 12'h0f0};
#337 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#337 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#338 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#338 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#339 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#339 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#340 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#340 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h055, 10'h000, 12'h105, 12'h0f0};
#340 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#341 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#341 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#341 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h055, 10'h000, 12'h105, 12'h0f0};
#342 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#342 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#343 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#343 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#344 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#344 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h056, 10'h000, 12'h106, 12'h0f0};
#344 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#345 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#345 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#345 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h056, 10'h000, 12'h106, 12'h0f0};
#346 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#346 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#347 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000a0, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000005, 32'h000000a0, 5'h09, 32'h000000a0, 32'h00004940, 32'h00000005, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#347 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a0, 32'h00000000, 32'h00000005};
#348 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000028, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000005, 32'h00000028, 5'h0a, 32'h00000028, 32'h000050c0, 32'h00000003, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#348 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h057, 10'h000, 12'h107, 12'h0f0};
#348 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000028, 32'h00000000, 32'h00000005};
#349 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000c8, 1'b0, 32'h00000000, 32'h00000028, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000a0, 32'h00000028, 32'h000000c8, 5'h09, 32'h000000c8, 32'h00004820, 32'h000000a0, 32'h00000028, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#349 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000c8, 32'h00000000, 32'h00000028};
#350 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000cd, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000c8, 32'h00000005, 32'h000000cd, 5'h09, 32'h000000cd, 32'h00004820, 32'h000000c8, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#350 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000cd, 32'h00000000, 32'h00000005};
#351 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000334, 1'b0, 32'h00000000, 32'h000000cd, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000cd, 32'h00000334, 5'h09, 32'h00000334, 32'h00004880, 32'h00000002, 32'h000000cd, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#351 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000334, 32'h00000000, 32'h000000cd};
#352 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020334, 1'b0, 32'h00000000, 32'h00000334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000334, 32'h10020334, 5'h08, 32'h10020334, 32'h00004020, 32'h10020000, 32'h00000334, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#352 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020334, 32'h00000000, 32'h00000334};
#352 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h058, 10'h000, 12'h108, 12'h0f0};
#353 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020334, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020334, 32'h00000002, 32'h10020334, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020334, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#353 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020334, 32'h00000000, 32'h00000002};
#353 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h058, 10'h000, 12'h108, 12'h0f0};
#354 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#354 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#354 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h058, 10'h000, 12'h108, 12'h0f0};
#355 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020334, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#355 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020334};
#356 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000334, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#356 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000334};
#356 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h059, 10'h000, 12'h109, 12'h0f0};
#357 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000028, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000028, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#357 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000028};
#358 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#358 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#359 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#359 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#360 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#360 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05a, 10'h000, 12'h10a, 12'h0f0};
#360 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#361 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#361 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#362 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#362 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#363 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#363 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#364 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#364 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05b, 10'h000, 12'h10b, 12'h0f0};
#364 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#365 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#365 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#365 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05b, 10'h000, 12'h10b, 12'h0f0};
#366 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#366 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#367 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#367 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#368 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#368 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05c, 10'h000, 12'h10c, 12'h0f0};
#368 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#369 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#369 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#369 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05c, 10'h000, 12'h10c, 12'h0f0};
#370 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#370 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#371 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000a0, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000005, 32'h000000a0, 5'h09, 32'h000000a0, 32'h00004940, 32'h00000005, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#371 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000a0, 32'h00000000, 32'h00000005};
#372 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000028, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000005, 32'h00000028, 5'h0a, 32'h00000028, 32'h000050c0, 32'h00000003, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#372 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05d, 10'h000, 12'h10d, 12'h0f0};
#372 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000028, 32'h00000000, 32'h00000005};
#373 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000c8, 1'b0, 32'h00000000, 32'h00000028, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000a0, 32'h00000028, 32'h000000c8, 5'h09, 32'h000000c8, 32'h00004820, 32'h000000a0, 32'h00000028, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#373 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000c8, 32'h00000000, 32'h00000028};
#374 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000cd, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000c8, 32'h00000005, 32'h000000cd, 5'h09, 32'h000000cd, 32'h00004820, 32'h000000c8, 32'h00000005, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#374 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000cd, 32'h00000000, 32'h00000005};
#375 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000334, 1'b0, 32'h00000000, 32'h000000cd, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000cd, 32'h00000334, 5'h09, 32'h00000334, 32'h00004880, 32'h00000002, 32'h000000cd, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#375 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000334, 32'h00000000, 32'h000000cd};
#376 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020334, 1'b0, 32'h00000002, 32'h00000334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000334, 32'h10020334, 5'h08, 32'h10020334, 32'h00004020, 32'h10020000, 32'h00000334, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#376 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020334, 32'h00000002, 32'h00000334};
#376 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05e, 10'h000, 12'h10e, 12'h0f0};
#377 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020334, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020334, 32'h00000003, 32'h10020334, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020334, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#377 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020334, 32'h00000002, 32'h00000003};
#377 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05e, 10'h000, 12'h10e, 12'h0f0};
#378 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#378 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#378 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05e, 10'h000, 12'h10e, 12'h0f0};
#379 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020334, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#379 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020334};
#380 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000334, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000334, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#380 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000334};
#380 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h005, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h05f, 10'h000, 12'h10f, 12'h0f0};
#381 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000028, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000028, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#381 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000028};
#382 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#382 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#383 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#383 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#384 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000006, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000006, 5'h05, 32'h00000006, 32'h00000001, 32'h00000005, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#384 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h060, 10'h000, 12'h200, 12'h00f};
#384 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000006, 32'h00000000, 32'h00000005};
#385 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000006, 1'b0, 32'h00000000, 32'h00000005, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000005, 32'h00000005, 32'h00000006, 5'h06, 32'h00000006, 32'h00000001, 32'h00000005, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#386 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000006, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000006, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#386 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#387 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#387 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#388 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#388 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h061, 10'h000, 12'h201, 12'h00f};
#388 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#389 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#389 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#390 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#390 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#391 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#391 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#391 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h061, 10'h000, 12'h201, 12'h00f};
#392 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#392 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#392 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h062, 10'h000, 12'h202, 12'h00f};
#393 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#393 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#394 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#394 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#395 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#395 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#395 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h062, 10'h000, 12'h202, 12'h00f};
#396 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#396 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h063, 10'h000, 12'h203, 12'h00f};
#396 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#397 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000c0, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000006, 32'h000000c0, 5'h09, 32'h000000c0, 32'h00004940, 32'h00000005, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#397 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000c0, 32'h00000000, 32'h00000006};
#398 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000030, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000006, 32'h00000030, 5'h0a, 32'h00000030, 32'h000050c0, 32'h00000003, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#398 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000030, 32'h00000000, 32'h00000006};
#399 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000f0, 1'b0, 32'h00000000, 32'h00000030, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000c0, 32'h00000030, 32'h000000f0, 5'h09, 32'h000000f0, 32'h00004820, 32'h000000c0, 32'h00000030, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#399 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000f0, 32'h00000000, 32'h00000030};
#400 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000f6, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000f0, 32'h00000006, 32'h000000f6, 5'h09, 32'h000000f6, 32'h00004820, 32'h000000f0, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#400 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000f6, 32'h00000000, 32'h00000006};
#400 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h064, 10'h000, 12'h204, 12'h00f};
#401 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000003d8, 1'b0, 32'h00000000, 32'h000000f6, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000f6, 32'h000003d8, 5'h09, 32'h000003d8, 32'h00004880, 32'h00000002, 32'h000000f6, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#401 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000003d8, 32'h00000000, 32'h000000f6};
#402 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100203d8, 1'b0, 32'h00000002, 32'h000003d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000003d8, 32'h100203d8, 5'h08, 32'h100203d8, 32'h00004020, 32'h10020000, 32'h000003d8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#402 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100203d8, 32'h00000002, 32'h000003d8};
#403 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100203d8, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100203d8, 32'h00000002, 32'h100203d8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100203d8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#403 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100203d8, 32'h00000002, 32'h00000002};
#403 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h064, 10'h000, 12'h204, 12'h00f};
#404 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#404 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h065, 10'h000, 12'h205, 12'h00f};
#404 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#405 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100203d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100203d8, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#405 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100203d8};
#406 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000003d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000003d8, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#406 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000003d8};
#407 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000030, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000030, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#407 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000030};
#408 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#408 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#408 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h066, 10'h000, 12'h206, 12'h00f};
#409 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#409 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#410 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#410 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#411 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#411 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#412 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#412 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h067, 10'h000, 12'h207, 12'h00f};
#412 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#413 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#413 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#414 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#414 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#415 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#415 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#415 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h067, 10'h000, 12'h207, 12'h00f};
#416 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#416 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#416 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h068, 10'h000, 12'h208, 12'h00f};
#417 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#417 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#418 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#418 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#419 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#419 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#419 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h068, 10'h000, 12'h208, 12'h00f};
#420 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#420 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h069, 10'h000, 12'h209, 12'h00f};
#420 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#421 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000c0, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000006, 32'h000000c0, 5'h09, 32'h000000c0, 32'h00004940, 32'h00000005, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#421 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000c0, 32'h00000000, 32'h00000006};
#422 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000030, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000006, 32'h00000030, 5'h0a, 32'h00000030, 32'h000050c0, 32'h00000003, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#422 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000030, 32'h00000000, 32'h00000006};
#423 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000000f0, 1'b0, 32'h00000000, 32'h00000030, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000c0, 32'h00000030, 32'h000000f0, 5'h09, 32'h000000f0, 32'h00004820, 32'h000000c0, 32'h00000030, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#423 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000f0, 32'h00000000, 32'h00000030};
#424 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000000f6, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000f0, 32'h00000006, 32'h000000f6, 5'h09, 32'h000000f6, 32'h00004820, 32'h000000f0, 32'h00000006, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#424 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000f6, 32'h00000000, 32'h00000006};
#424 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06a, 10'h000, 12'h20a, 12'h00f};
#425 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000003d8, 1'b0, 32'h00000000, 32'h000000f6, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000f6, 32'h000003d8, 5'h09, 32'h000003d8, 32'h00004880, 32'h00000002, 32'h000000f6, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#425 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000003d8, 32'h00000000, 32'h000000f6};
#426 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100203d8, 1'b0, 32'h00000002, 32'h000003d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000003d8, 32'h100203d8, 5'h08, 32'h100203d8, 32'h00004020, 32'h10020000, 32'h000003d8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#426 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100203d8, 32'h00000002, 32'h000003d8};
#427 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100203d8, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100203d8, 32'h00000003, 32'h100203d8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100203d8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#427 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100203d8, 32'h00000002, 32'h00000003};
#427 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06a, 10'h000, 12'h20a, 12'h00f};
#428 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#428 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#428 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06b, 10'h000, 12'h20b, 12'h00f};
#429 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100203d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100203d8, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#429 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100203d8};
#430 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000003d8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000003d8, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#430 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000003d8};
#431 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000030, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000030, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#431 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000030};
#432 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#432 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#432 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06c, 10'h000, 12'h20c, 12'h00f};
#433 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#433 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#434 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000007, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000006, 32'h00000006, 32'h00000007, 5'h05, 32'h00000007, 32'h00000001, 32'h00000006, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#434 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000000, 32'h00000007, 32'h00000000, 32'h00000006};
#435 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000007, 1'b0, 32'h00000000, 32'h00000006, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000006, 32'h00000006, 32'h00000007, 5'h06, 32'h00000007, 32'h00000001, 32'h00000006, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#436 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000007, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000007, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#436 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#436 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06d, 10'h000, 12'h20d, 12'h00f};
#437 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#437 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#438 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#438 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#439 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#439 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#440 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#440 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06e, 10'h000, 12'h20e, 12'h00f};
#440 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#441 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#441 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#441 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06e, 10'h000, 12'h20e, 12'h00f};
#442 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#442 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#443 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#443 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#444 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#444 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06f, 10'h000, 12'h20f, 12'h00f};
#444 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#445 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#445 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#445 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h006, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h06f, 10'h000, 12'h20f, 12'h00f};
#446 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#446 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#447 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000e0, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000007, 32'h000000e0, 5'h09, 32'h000000e0, 32'h00004940, 32'h00000005, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#447 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000e0, 32'h00000000, 32'h00000007};
#448 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000038, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000007, 32'h00000038, 5'h0a, 32'h00000038, 32'h000050c0, 32'h00000003, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#448 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h070, 10'h000, 12'h200, 12'h00f};
#448 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000038, 32'h00000000, 32'h00000007};
#449 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000118, 1'b0, 32'h00000000, 32'h00000038, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000e0, 32'h00000038, 32'h00000118, 5'h09, 32'h00000118, 32'h00004820, 32'h000000e0, 32'h00000038, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#449 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000118, 32'h00000000, 32'h00000038};
#450 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000011f, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000118, 32'h00000007, 32'h0000011f, 5'h09, 32'h0000011f, 32'h00004820, 32'h00000118, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#450 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000011f, 32'h00000000, 32'h00000007};
#451 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000047c, 1'b0, 32'h00000000, 32'h0000011f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000011f, 32'h0000047c, 5'h09, 32'h0000047c, 32'h00004880, 32'h00000002, 32'h0000011f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#451 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000047c, 32'h00000000, 32'h0000011f};
#452 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002047c, 1'b0, 32'h00000003, 32'h0000047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000047c, 32'h1002047c, 5'h08, 32'h1002047c, 32'h00004020, 32'h10020000, 32'h0000047c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#452 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002047c, 32'h00000003, 32'h0000047c};
#452 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h071, 10'h000, 12'h201, 12'h00f};
#453 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002047c, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002047c, 32'h00000002, 32'h1002047c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002047c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#453 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002047c, 32'h00000003, 32'h00000002};
#453 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h071, 10'h000, 12'h201, 12'h00f};
#454 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#454 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#454 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h071, 10'h000, 12'h201, 12'h00f};
#455 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002047c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#455 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002047c};
#456 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000047c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#456 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000047c};
#456 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h072, 10'h000, 12'h202, 12'h00f};
#457 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000038, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000038, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#457 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000038};
#458 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#458 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#459 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#459 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#460 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#460 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h073, 10'h000, 12'h203, 12'h00f};
#460 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#461 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#461 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#462 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#462 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#463 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#463 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#464 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#464 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h074, 10'h000, 12'h204, 12'h00f};
#464 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#465 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#465 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#465 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h074, 10'h000, 12'h204, 12'h00f};
#466 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#466 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#467 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#467 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#468 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#468 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h075, 10'h000, 12'h205, 12'h00f};
#468 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#469 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#469 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#469 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h075, 10'h000, 12'h205, 12'h00f};
#470 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#470 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#471 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000000e0, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000007, 32'h000000e0, 5'h09, 32'h000000e0, 32'h00004940, 32'h00000005, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#471 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000000e0, 32'h00000000, 32'h00000007};
#472 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000038, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000007, 32'h00000038, 5'h0a, 32'h00000038, 32'h000050c0, 32'h00000003, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#472 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h076, 10'h000, 12'h206, 12'h00f};
#472 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000038, 32'h00000000, 32'h00000007};
#473 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000118, 1'b0, 32'h00000000, 32'h00000038, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000000e0, 32'h00000038, 32'h00000118, 5'h09, 32'h00000118, 32'h00004820, 32'h000000e0, 32'h00000038, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#473 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000118, 32'h00000000, 32'h00000038};
#474 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000011f, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000118, 32'h00000007, 32'h0000011f, 5'h09, 32'h0000011f, 32'h00004820, 32'h00000118, 32'h00000007, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#474 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000011f, 32'h00000000, 32'h00000007};
#475 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000047c, 1'b0, 32'h00000000, 32'h0000011f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000011f, 32'h0000047c, 5'h09, 32'h0000047c, 32'h00004880, 32'h00000002, 32'h0000011f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#475 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000047c, 32'h00000000, 32'h0000011f};
#476 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002047c, 1'b0, 32'h00000002, 32'h0000047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000047c, 32'h1002047c, 5'h08, 32'h1002047c, 32'h00004020, 32'h10020000, 32'h0000047c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#476 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002047c, 32'h00000002, 32'h0000047c};
#476 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h077, 10'h000, 12'h207, 12'h00f};
#477 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002047c, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002047c, 32'h00000003, 32'h1002047c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002047c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#477 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002047c, 32'h00000002, 32'h00000003};
#477 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h077, 10'h000, 12'h207, 12'h00f};
#478 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#478 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#478 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h077, 10'h000, 12'h207, 12'h00f};
#479 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002047c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#479 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002047c};
#480 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000047c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000047c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#480 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000047c};
#480 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h078, 10'h000, 12'h208, 12'h00f};
#481 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000038, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000038, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#481 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000038};
#482 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#482 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#483 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#483 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#484 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000008, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000007, 32'h00000007, 32'h00000008, 5'h05, 32'h00000008, 32'h00000001, 32'h00000007, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#484 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h079, 10'h000, 12'h209, 12'h00f};
#484 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000008, 32'h00000000, 32'h00000007};
#485 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000008, 1'b0, 32'h00000000, 32'h00000007, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000007, 32'h00000007, 32'h00000008, 5'h06, 32'h00000008, 32'h00000001, 32'h00000007, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#486 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000008, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000008, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#486 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#487 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#487 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#488 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#488 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07a, 10'h000, 12'h20a, 12'h00f};
#488 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#489 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#489 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#490 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#490 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#491 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#491 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#491 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07a, 10'h000, 12'h20a, 12'h00f};
#492 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#492 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#492 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07b, 10'h000, 12'h20b, 12'h00f};
#493 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#493 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#494 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#494 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#495 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#495 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#495 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07b, 10'h000, 12'h20b, 12'h00f};
#496 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#496 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07c, 10'h000, 12'h20c, 12'h00f};
#496 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#497 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000100, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000100, 5'h09, 32'h00000100, 32'h00004940, 32'h00000005, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#497 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000100, 32'h00000000, 32'h00000008};
#498 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000040, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000040, 5'h0a, 32'h00000040, 32'h000050c0, 32'h00000003, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#498 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000040, 32'h00000000, 32'h00000008};
#499 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000140, 1'b0, 32'h00000000, 32'h00000040, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000100, 32'h00000040, 32'h00000140, 5'h09, 32'h00000140, 32'h00004820, 32'h00000100, 32'h00000040, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#499 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000140, 32'h00000000, 32'h00000040};
#500 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000148, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000140, 32'h00000008, 32'h00000148, 5'h09, 32'h00000148, 32'h00004820, 32'h00000140, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#500 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000148, 32'h00000000, 32'h00000008};
#500 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07d, 10'h000, 12'h20d, 12'h00f};
#501 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000520, 1'b0, 32'h00000000, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000148, 32'h00000520, 5'h09, 32'h00000520, 32'h00004880, 32'h00000002, 32'h00000148, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#501 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000520, 32'h00000000, 32'h00000148};
#502 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020520, 1'b0, 32'h00000001, 32'h00000520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000520, 32'h10020520, 5'h08, 32'h10020520, 32'h00004020, 32'h10020000, 32'h00000520, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#502 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020520, 32'h00000001, 32'h00000520};
#503 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020520, 1'b1, 32'h00000001, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020520, 32'h00000002, 32'h10020520, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020520, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#503 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020520, 32'h00000001, 32'h00000002};
#503 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07d, 10'h000, 12'h20d, 12'h00f};
#504 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#504 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#504 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07e, 10'h000, 12'h20e, 12'h00f};
#505 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020520, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#505 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020520};
#506 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000520, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#506 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000520};
#507 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000040, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000040, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#507 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000040};
#508 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#508 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#508 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h007, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h07f, 10'h000, 12'h20f, 12'h00f};
#509 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#509 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#510 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#510 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#511 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#511 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#512 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#512 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h080, 10'h000, 12'h200, 12'h00f};
#512 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#513 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#513 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#514 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#514 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#515 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#515 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#515 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h080, 10'h000, 12'h200, 12'h00f};
#516 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#516 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#516 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h081, 10'h000, 12'h201, 12'h00f};
#517 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#517 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#518 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#518 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#519 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#519 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#519 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h081, 10'h000, 12'h201, 12'h00f};
#520 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#520 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h082, 10'h000, 12'h202, 12'h00f};
#520 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#521 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000100, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000100, 5'h09, 32'h00000100, 32'h00004940, 32'h00000005, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#521 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000100, 32'h00000000, 32'h00000008};
#522 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000040, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000040, 5'h0a, 32'h00000040, 32'h000050c0, 32'h00000003, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#522 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000040, 32'h00000000, 32'h00000008};
#523 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000140, 1'b0, 32'h00000000, 32'h00000040, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000100, 32'h00000040, 32'h00000140, 5'h09, 32'h00000140, 32'h00004820, 32'h00000100, 32'h00000040, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#523 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000140, 32'h00000000, 32'h00000040};
#524 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000148, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000140, 32'h00000008, 32'h00000148, 5'h09, 32'h00000148, 32'h00004820, 32'h00000140, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#524 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000148, 32'h00000000, 32'h00000008};
#524 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h083, 10'h000, 12'h203, 12'h00f};
#525 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000520, 1'b0, 32'h00000000, 32'h00000148, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000148, 32'h00000520, 5'h09, 32'h00000520, 32'h00004880, 32'h00000002, 32'h00000148, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#525 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000520, 32'h00000000, 32'h00000148};
#526 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020520, 1'b0, 32'h00000002, 32'h00000520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000520, 32'h10020520, 5'h08, 32'h10020520, 32'h00004020, 32'h10020000, 32'h00000520, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#526 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020520, 32'h00000002, 32'h00000520};
#527 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020520, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020520, 32'h00000003, 32'h10020520, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020520, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#527 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020520, 32'h00000002, 32'h00000003};
#527 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h083, 10'h000, 12'h203, 12'h00f};
#528 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#528 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#528 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h084, 10'h000, 12'h204, 12'h00f};
#529 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020520, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#529 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020520};
#530 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000520, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000520, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#530 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000520};
#531 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000040, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000040, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#531 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000040};
#532 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#532 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#532 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h085, 10'h000, 12'h205, 12'h00f};
#533 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#533 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#534 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000009, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h00000009, 5'h05, 32'h00000009, 32'h00000001, 32'h00000008, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#534 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000009, 32'h00000000, 32'h00000008};
#535 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000009, 1'b0, 32'h00000000, 32'h00000008, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h00000009, 5'h06, 32'h00000009, 32'h00000001, 32'h00000008, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#536 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000009, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000009, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#536 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#536 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h086, 10'h000, 12'h206, 12'h00f};
#537 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#537 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#538 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#538 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#539 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#539 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#540 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#540 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h087, 10'h000, 12'h207, 12'h00f};
#540 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#541 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#541 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#541 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h087, 10'h000, 12'h207, 12'h00f};
#542 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#542 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#543 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#543 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#544 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#544 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h088, 10'h000, 12'h208, 12'h00f};
#544 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#545 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#545 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#545 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h088, 10'h000, 12'h208, 12'h00f};
#546 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#546 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#547 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000120, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000009, 32'h00000120, 5'h09, 32'h00000120, 32'h00004940, 32'h00000005, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#547 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000120, 32'h00000000, 32'h00000009};
#548 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000048, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000009, 32'h00000048, 5'h0a, 32'h00000048, 32'h000050c0, 32'h00000003, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#548 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h089, 10'h000, 12'h209, 12'h00f};
#548 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000048, 32'h00000000, 32'h00000009};
#549 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000168, 1'b0, 32'h00000000, 32'h00000048, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000120, 32'h00000048, 32'h00000168, 5'h09, 32'h00000168, 32'h00004820, 32'h00000120, 32'h00000048, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#549 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000168, 32'h00000000, 32'h00000048};
#550 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000171, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000168, 32'h00000009, 32'h00000171, 5'h09, 32'h00000171, 32'h00004820, 32'h00000168, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#550 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000171, 32'h00000000, 32'h00000009};
#551 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000005c4, 1'b0, 32'h00000000, 32'h00000171, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000171, 32'h000005c4, 5'h09, 32'h000005c4, 32'h00004880, 32'h00000002, 32'h00000171, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#551 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000005c4, 32'h00000000, 32'h00000171};
#552 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100205c4, 1'b0, 32'h00000003, 32'h000005c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000005c4, 32'h100205c4, 5'h08, 32'h100205c4, 32'h00004020, 32'h10020000, 32'h000005c4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#552 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100205c4, 32'h00000003, 32'h000005c4};
#552 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08a, 10'h000, 12'h20a, 12'h00f};
#553 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100205c4, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100205c4, 32'h00000002, 32'h100205c4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100205c4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#553 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100205c4, 32'h00000003, 32'h00000002};
#553 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08a, 10'h000, 12'h20a, 12'h00f};
#554 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#554 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#554 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08a, 10'h000, 12'h20a, 12'h00f};
#555 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100205c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100205c4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#555 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100205c4};
#556 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000005c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000005c4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#556 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000005c4};
#556 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08b, 10'h000, 12'h20b, 12'h00f};
#557 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000048, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000048, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#557 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000048};
#558 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#558 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#559 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#559 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#560 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#560 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08c, 10'h000, 12'h20c, 12'h00f};
#560 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#561 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#561 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#562 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#562 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#563 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#563 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#564 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#564 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08d, 10'h000, 12'h20d, 12'h00f};
#564 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#565 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#565 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#565 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08d, 10'h000, 12'h20d, 12'h00f};
#566 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#566 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#567 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#567 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#568 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#568 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08e, 10'h000, 12'h20e, 12'h00f};
#568 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#569 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#569 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#569 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08e, 10'h000, 12'h20e, 12'h00f};
#570 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#570 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#571 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000120, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000009, 32'h00000120, 5'h09, 32'h00000120, 32'h00004940, 32'h00000005, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#571 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000120, 32'h00000000, 32'h00000009};
#572 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000048, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000009, 32'h00000048, 5'h0a, 32'h00000048, 32'h000050c0, 32'h00000003, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#572 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h008, 4'h2, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'h0, 4'hf, 10'h08f, 10'h000, 12'h20f, 12'h00f};
#572 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000048, 32'h00000000, 32'h00000009};
#573 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000168, 1'b0, 32'h00000000, 32'h00000048, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000120, 32'h00000048, 32'h00000168, 5'h09, 32'h00000168, 32'h00004820, 32'h00000120, 32'h00000048, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#573 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000168, 32'h00000000, 32'h00000048};
#574 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000171, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000168, 32'h00000009, 32'h00000171, 5'h09, 32'h00000171, 32'h00004820, 32'h00000168, 32'h00000009, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#574 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000171, 32'h00000000, 32'h00000009};
#575 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000005c4, 1'b0, 32'h00000000, 32'h00000171, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000171, 32'h000005c4, 5'h09, 32'h000005c4, 32'h00004880, 32'h00000002, 32'h00000171, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#575 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000005c4, 32'h00000000, 32'h00000171};
#576 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100205c4, 1'b0, 32'h00000002, 32'h000005c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000005c4, 32'h100205c4, 5'h08, 32'h100205c4, 32'h00004020, 32'h10020000, 32'h000005c4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#576 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100205c4, 32'h00000002, 32'h000005c4};
#576 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h090, 10'h000, 12'h300, 12'hfff};
#577 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100205c4, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100205c4, 32'h00000003, 32'h100205c4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100205c4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#577 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100205c4, 32'h00000002, 32'h00000003};
#577 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h090, 10'h000, 12'h300, 12'hfff};
#578 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#578 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#578 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h090, 10'h000, 12'h300, 12'hfff};
#579 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100205c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100205c4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#579 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100205c4};
#580 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000005c4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000005c4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#580 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000005c4};
#580 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h091, 10'h000, 12'h301, 12'hfff};
#581 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000048, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000048, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#581 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000048};
#582 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#582 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#583 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#583 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#584 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000a, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000009, 32'h00000009, 32'h0000000a, 5'h05, 32'h0000000a, 32'h00000001, 32'h00000009, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#584 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h092, 10'h000, 12'h302, 12'hfff};
#584 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000a, 32'h00000000, 32'h00000009};
#585 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000a, 1'b0, 32'h00000000, 32'h00000009, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000009, 32'h00000009, 32'h0000000a, 5'h06, 32'h0000000a, 32'h00000001, 32'h00000009, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#586 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000a, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000a, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#586 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#587 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#587 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#588 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#588 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h093, 10'h000, 12'h303, 12'hfff};
#588 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#589 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#589 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#590 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#590 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#591 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#591 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#591 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h093, 10'h000, 12'h303, 12'hfff};
#592 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#592 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#592 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h094, 10'h000, 12'h304, 12'hfff};
#593 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#593 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#594 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#594 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#595 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#595 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#595 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h094, 10'h000, 12'h304, 12'hfff};
#596 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#596 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h095, 10'h000, 12'h305, 12'hfff};
#596 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#597 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000140, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000140, 5'h09, 32'h00000140, 32'h00004940, 32'h00000005, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#597 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000140, 32'h00000000, 32'h0000000a};
#598 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000050, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000050, 5'h0a, 32'h00000050, 32'h000050c0, 32'h00000003, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#598 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000050, 32'h00000000, 32'h0000000a};
#599 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000190, 1'b0, 32'h00000000, 32'h00000050, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000140, 32'h00000050, 32'h00000190, 5'h09, 32'h00000190, 32'h00004820, 32'h00000140, 32'h00000050, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#599 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000190, 32'h00000000, 32'h00000050};
#600 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000019a, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000190, 32'h0000000a, 32'h0000019a, 5'h09, 32'h0000019a, 32'h00004820, 32'h00000190, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#600 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000019a, 32'h00000000, 32'h0000000a};
#600 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h096, 10'h000, 12'h306, 12'hfff};
#601 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000668, 1'b0, 32'h00000000, 32'h0000019a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000019a, 32'h00000668, 5'h09, 32'h00000668, 32'h00004880, 32'h00000002, 32'h0000019a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#601 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000668, 32'h00000000, 32'h0000019a};
#602 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020668, 1'b0, 32'h00000000, 32'h00000668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000668, 32'h10020668, 5'h08, 32'h10020668, 32'h00004020, 32'h10020000, 32'h00000668, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#602 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020668, 32'h00000000, 32'h00000668};
#603 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020668, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020668, 32'h00000002, 32'h10020668, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020668, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#603 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020668, 32'h00000000, 32'h00000002};
#603 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h096, 10'h000, 12'h306, 12'hfff};
#604 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#604 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#604 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h097, 10'h000, 12'h307, 12'hfff};
#605 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020668, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#605 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020668};
#606 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000668, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#606 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000668};
#607 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000050, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000050, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#607 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000050};
#608 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#608 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#608 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h098, 10'h000, 12'h308, 12'hfff};
#609 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#609 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#610 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#610 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#611 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#611 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#612 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#612 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h099, 10'h000, 12'h309, 12'hfff};
#612 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#613 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#613 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#614 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#614 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#615 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#615 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#615 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h099, 10'h000, 12'h309, 12'hfff};
#616 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#616 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#616 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09a, 10'h000, 12'h30a, 12'hfff};
#617 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#617 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#618 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#618 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#619 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#619 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#619 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09a, 10'h000, 12'h30a, 12'hfff};
#620 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#620 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09b, 10'h000, 12'h30b, 12'hfff};
#620 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#621 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000140, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000140, 5'h09, 32'h00000140, 32'h00004940, 32'h00000005, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#621 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000140, 32'h00000000, 32'h0000000a};
#622 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000050, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000050, 5'h0a, 32'h00000050, 32'h000050c0, 32'h00000003, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#622 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000050, 32'h00000000, 32'h0000000a};
#623 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000190, 1'b0, 32'h00000000, 32'h00000050, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000140, 32'h00000050, 32'h00000190, 5'h09, 32'h00000190, 32'h00004820, 32'h00000140, 32'h00000050, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#623 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000190, 32'h00000000, 32'h00000050};
#624 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000019a, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000190, 32'h0000000a, 32'h0000019a, 5'h09, 32'h0000019a, 32'h00004820, 32'h00000190, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#624 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000019a, 32'h00000000, 32'h0000000a};
#624 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09c, 10'h000, 12'h30c, 12'hfff};
#625 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000668, 1'b0, 32'h00000000, 32'h0000019a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000019a, 32'h00000668, 5'h09, 32'h00000668, 32'h00004880, 32'h00000002, 32'h0000019a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#625 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000668, 32'h00000000, 32'h0000019a};
#626 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020668, 1'b0, 32'h00000002, 32'h00000668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000668, 32'h10020668, 5'h08, 32'h10020668, 32'h00004020, 32'h10020000, 32'h00000668, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#626 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020668, 32'h00000002, 32'h00000668};
#627 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020668, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020668, 32'h00000003, 32'h10020668, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020668, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#627 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020668, 32'h00000002, 32'h00000003};
#627 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09c, 10'h000, 12'h30c, 12'hfff};
#628 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#628 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#628 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09d, 10'h000, 12'h30d, 12'hfff};
#629 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020668, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#629 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020668};
#630 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000668, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000668, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#630 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000668};
#631 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000050, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000050, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#631 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000050};
#632 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#632 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#632 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09e, 10'h000, 12'h30e, 12'hfff};
#633 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#633 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#634 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000b, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000a, 32'h0000000a, 32'h0000000b, 5'h05, 32'h0000000b, 32'h00000001, 32'h0000000a, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#634 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000b, 32'h00000000, 32'h0000000a};
#635 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000b, 1'b0, 32'h00000000, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000a, 32'h0000000a, 32'h0000000b, 5'h06, 32'h0000000b, 32'h00000001, 32'h0000000a, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#636 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000b, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000b, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#636 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#636 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h009, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h09f, 10'h000, 12'h30f, 12'hfff};
#637 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#637 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#638 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#638 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#639 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#639 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#640 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#640 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a0, 10'h000, 12'h300, 12'hfff};
#640 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#641 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#641 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#641 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a0, 10'h000, 12'h300, 12'hfff};
#642 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#642 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#643 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#643 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#644 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#644 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a1, 10'h000, 12'h301, 12'hfff};
#644 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#645 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#645 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#645 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a1, 10'h000, 12'h301, 12'hfff};
#646 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#646 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#647 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000160, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000160, 5'h09, 32'h00000160, 32'h00004940, 32'h00000005, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#647 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000160, 32'h00000000, 32'h0000000b};
#648 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000058, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000058, 5'h0a, 32'h00000058, 32'h000050c0, 32'h00000003, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#648 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a2, 10'h000, 12'h302, 12'hfff};
#648 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000058, 32'h00000000, 32'h0000000b};
#649 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000001b8, 1'b0, 32'h00000000, 32'h00000058, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000160, 32'h00000058, 32'h000001b8, 5'h09, 32'h000001b8, 32'h00004820, 32'h00000160, 32'h00000058, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#649 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001b8, 32'h00000000, 32'h00000058};
#650 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000001c3, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001b8, 32'h0000000b, 32'h000001c3, 5'h09, 32'h000001c3, 32'h00004820, 32'h000001b8, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#650 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001c3, 32'h00000000, 32'h0000000b};
#651 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000070c, 1'b0, 32'h00000000, 32'h000001c3, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001c3, 32'h0000070c, 5'h09, 32'h0000070c, 32'h00004880, 32'h00000002, 32'h000001c3, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#651 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000070c, 32'h00000000, 32'h000001c3};
#652 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002070c, 1'b0, 32'h00000002, 32'h0000070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000070c, 32'h1002070c, 5'h08, 32'h1002070c, 32'h00004020, 32'h10020000, 32'h0000070c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#652 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002070c, 32'h00000002, 32'h0000070c};
#652 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a3, 10'h000, 12'h303, 12'hfff};
#653 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002070c, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002070c, 32'h00000002, 32'h1002070c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002070c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#653 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002070c, 32'h00000002, 32'h00000002};
#653 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a3, 10'h000, 12'h303, 12'hfff};
#654 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#654 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#654 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a3, 10'h000, 12'h303, 12'hfff};
#655 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002070c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#655 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002070c};
#656 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000070c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#656 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000070c};
#656 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a4, 10'h000, 12'h304, 12'hfff};
#657 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000058, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000058, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#657 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000058};
#658 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#658 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#659 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#659 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#660 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#660 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a5, 10'h000, 12'h305, 12'hfff};
#660 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#661 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#661 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#662 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#662 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#663 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#663 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#664 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#664 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a6, 10'h000, 12'h306, 12'hfff};
#664 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#665 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#665 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#665 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a6, 10'h000, 12'h306, 12'hfff};
#666 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#666 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#667 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#667 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#668 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#668 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a7, 10'h000, 12'h307, 12'hfff};
#668 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#669 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#669 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#669 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a7, 10'h000, 12'h307, 12'hfff};
#670 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#670 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#671 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000160, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000160, 5'h09, 32'h00000160, 32'h00004940, 32'h00000005, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#671 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000160, 32'h00000000, 32'h0000000b};
#672 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000058, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000058, 5'h0a, 32'h00000058, 32'h000050c0, 32'h00000003, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#672 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a8, 10'h000, 12'h308, 12'hfff};
#672 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000058, 32'h00000000, 32'h0000000b};
#673 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000001b8, 1'b0, 32'h00000000, 32'h00000058, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000160, 32'h00000058, 32'h000001b8, 5'h09, 32'h000001b8, 32'h00004820, 32'h00000160, 32'h00000058, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#673 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001b8, 32'h00000000, 32'h00000058};
#674 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000001c3, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001b8, 32'h0000000b, 32'h000001c3, 5'h09, 32'h000001c3, 32'h00004820, 32'h000001b8, 32'h0000000b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#674 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001c3, 32'h00000000, 32'h0000000b};
#675 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000070c, 1'b0, 32'h00000000, 32'h000001c3, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001c3, 32'h0000070c, 5'h09, 32'h0000070c, 32'h00004880, 32'h00000002, 32'h000001c3, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#675 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000070c, 32'h00000000, 32'h000001c3};
#676 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002070c, 1'b0, 32'h00000002, 32'h0000070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000070c, 32'h1002070c, 5'h08, 32'h1002070c, 32'h00004020, 32'h10020000, 32'h0000070c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#676 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002070c, 32'h00000002, 32'h0000070c};
#676 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a9, 10'h000, 12'h309, 12'hfff};
#677 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002070c, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002070c, 32'h00000003, 32'h1002070c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002070c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#677 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002070c, 32'h00000002, 32'h00000003};
#677 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a9, 10'h000, 12'h309, 12'hfff};
#678 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#678 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#678 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0a9, 10'h000, 12'h309, 12'hfff};
#679 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002070c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#679 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002070c};
#680 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000070c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000070c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#680 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000070c};
#680 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0aa, 10'h000, 12'h30a, 12'hfff};
#681 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000058, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000058, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#681 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000058};
#682 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#682 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#683 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#683 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#684 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000c, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000b, 32'h0000000b, 32'h0000000c, 5'h05, 32'h0000000c, 32'h00000001, 32'h0000000b, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#684 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ab, 10'h000, 12'h30b, 12'hfff};
#684 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000c, 32'h00000000, 32'h0000000b};
#685 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000c, 1'b0, 32'h00000000, 32'h0000000b, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000b, 32'h0000000b, 32'h0000000c, 5'h06, 32'h0000000c, 32'h00000001, 32'h0000000b, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#686 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000c, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000c, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#686 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#687 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#687 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#688 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#688 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ac, 10'h000, 12'h30c, 12'hfff};
#688 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#689 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#689 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#690 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#690 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#691 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#691 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#691 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ac, 10'h000, 12'h30c, 12'hfff};
#692 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#692 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#692 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ad, 10'h000, 12'h30d, 12'hfff};
#693 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#693 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#694 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#694 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#695 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#695 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#695 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ad, 10'h000, 12'h30d, 12'hfff};
#696 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#696 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ae, 10'h000, 12'h30e, 12'hfff};
#696 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#697 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000180, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000180, 5'h09, 32'h00000180, 32'h00004940, 32'h00000005, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#697 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000180, 32'h00000000, 32'h0000000c};
#698 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000060, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000060, 5'h0a, 32'h00000060, 32'h000050c0, 32'h00000003, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#698 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000060, 32'h00000000, 32'h0000000c};
#699 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000001e0, 1'b0, 32'h00000000, 32'h00000060, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000180, 32'h00000060, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004820, 32'h00000180, 32'h00000060, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#699 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001e0, 32'h00000000, 32'h00000060};
#700 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000001ec, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h0000000c, 32'h000001ec, 5'h09, 32'h000001ec, 32'h00004820, 32'h000001e0, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#700 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001ec, 32'h00000000, 32'h0000000c};
#700 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0af, 10'h000, 12'h30f, 12'hfff};
#701 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000007b0, 1'b0, 32'h00000000, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001ec, 32'h000007b0, 5'h09, 32'h000007b0, 32'h00004880, 32'h00000002, 32'h000001ec, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#701 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000007b0, 32'h00000000, 32'h000001ec};
#702 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100207b0, 1'b0, 32'h00000000, 32'h000007b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000007b0, 32'h100207b0, 5'h08, 32'h100207b0, 32'h00004020, 32'h10020000, 32'h000007b0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#702 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100207b0, 32'h00000000, 32'h000007b0};
#703 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100207b0, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100207b0, 32'h00000002, 32'h100207b0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100207b0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#703 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100207b0, 32'h00000000, 32'h00000002};
#703 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00a, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0af, 10'h000, 12'h30f, 12'hfff};
#704 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#704 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#704 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b0, 10'h000, 12'h300, 12'hfff};
#705 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100207b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100207b0, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#705 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100207b0};
#706 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000007b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000007b0, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#706 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000007b0};
#707 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000060, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000060, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#707 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000060};
#708 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#708 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#708 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b1, 10'h000, 12'h301, 12'hfff};
#709 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#709 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#710 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#710 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#711 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#711 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#712 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#712 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b2, 10'h000, 12'h302, 12'hfff};
#712 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#713 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#713 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#714 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#714 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#715 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#715 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#715 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b2, 10'h000, 12'h302, 12'hfff};
#716 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#716 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#716 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b3, 10'h000, 12'h303, 12'hfff};
#717 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#717 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#718 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#718 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#719 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#719 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#719 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b3, 10'h000, 12'h303, 12'hfff};
#720 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#720 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b4, 10'h000, 12'h304, 12'hfff};
#720 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#721 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000180, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000180, 5'h09, 32'h00000180, 32'h00004940, 32'h00000005, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#721 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000180, 32'h00000000, 32'h0000000c};
#722 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000060, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000060, 5'h0a, 32'h00000060, 32'h000050c0, 32'h00000003, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#722 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000060, 32'h00000000, 32'h0000000c};
#723 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000001e0, 1'b0, 32'h00000000, 32'h00000060, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000180, 32'h00000060, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004820, 32'h00000180, 32'h00000060, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#723 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001e0, 32'h00000000, 32'h00000060};
#724 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000001ec, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h0000000c, 32'h000001ec, 5'h09, 32'h000001ec, 32'h00004820, 32'h000001e0, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#724 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001ec, 32'h00000000, 32'h0000000c};
#724 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b5, 10'h000, 12'h305, 12'hfff};
#725 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000007b0, 1'b0, 32'h00000000, 32'h000001ec, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001ec, 32'h000007b0, 5'h09, 32'h000007b0, 32'h00004880, 32'h00000002, 32'h000001ec, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#725 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000007b0, 32'h00000000, 32'h000001ec};
#726 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100207b0, 1'b0, 32'h00000002, 32'h000007b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000007b0, 32'h100207b0, 5'h08, 32'h100207b0, 32'h00004020, 32'h10020000, 32'h000007b0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#726 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100207b0, 32'h00000002, 32'h000007b0};
#727 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100207b0, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100207b0, 32'h00000003, 32'h100207b0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100207b0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#727 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100207b0, 32'h00000002, 32'h00000003};
#727 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b5, 10'h000, 12'h305, 12'hfff};
#728 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#728 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#728 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b6, 10'h000, 12'h306, 12'hfff};
#729 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100207b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100207b0, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#729 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100207b0};
#730 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000007b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000007b0, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#730 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000007b0};
#731 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000060, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000060, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#731 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000060};
#732 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#732 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#732 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b7, 10'h000, 12'h307, 12'hfff};
#733 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#733 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#734 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000d, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000c, 32'h0000000c, 32'h0000000d, 5'h05, 32'h0000000d, 32'h00000001, 32'h0000000c, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#734 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000d, 32'h00000000, 32'h0000000c};
#735 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000d, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000c, 32'h0000000c, 32'h0000000d, 5'h06, 32'h0000000d, 32'h00000001, 32'h0000000c, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#736 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000d, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000d, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#736 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#736 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b8, 10'h000, 12'h308, 12'hfff};
#737 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#737 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#738 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#738 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#739 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#739 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#740 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#740 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b9, 10'h000, 12'h309, 12'hfff};
#740 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#741 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#741 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#741 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0b9, 10'h000, 12'h309, 12'hfff};
#742 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#742 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#743 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#743 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#744 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#744 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ba, 10'h000, 12'h30a, 12'hfff};
#744 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#745 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#745 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#745 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ba, 10'h000, 12'h30a, 12'hfff};
#746 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#746 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#747 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001a0, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h000001a0, 5'h09, 32'h000001a0, 32'h00004940, 32'h00000005, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#747 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001a0, 32'h00000000, 32'h0000000d};
#748 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000068, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000068, 5'h0a, 32'h00000068, 32'h000050c0, 32'h00000003, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#748 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bb, 10'h000, 12'h30b, 12'hfff};
#748 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000068, 32'h00000000, 32'h0000000d};
#749 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000208, 1'b0, 32'h00000000, 32'h00000068, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001a0, 32'h00000068, 32'h00000208, 5'h09, 32'h00000208, 32'h00004820, 32'h000001a0, 32'h00000068, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#749 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000208, 32'h00000000, 32'h00000068};
#750 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000215, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000208, 32'h0000000d, 32'h00000215, 5'h09, 32'h00000215, 32'h00004820, 32'h00000208, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#750 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000215, 32'h00000000, 32'h0000000d};
#751 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000854, 1'b0, 32'h00000000, 32'h00000215, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000215, 32'h00000854, 5'h09, 32'h00000854, 32'h00004880, 32'h00000002, 32'h00000215, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#751 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000854, 32'h00000000, 32'h00000215};
#752 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020854, 1'b0, 32'h00000001, 32'h00000854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000854, 32'h10020854, 5'h08, 32'h10020854, 32'h00004020, 32'h10020000, 32'h00000854, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#752 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020854, 32'h00000001, 32'h00000854};
#752 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bc, 10'h000, 12'h30c, 12'hfff};
#753 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020854, 1'b1, 32'h00000001, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020854, 32'h00000002, 32'h10020854, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020854, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#753 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020854, 32'h00000001, 32'h00000002};
#753 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bc, 10'h000, 12'h30c, 12'hfff};
#754 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#754 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#754 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bc, 10'h000, 12'h30c, 12'hfff};
#755 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020854, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#755 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020854};
#756 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000854, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#756 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000854};
#756 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bd, 10'h000, 12'h30d, 12'hfff};
#757 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000068, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000068, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#757 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000068};
#758 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#758 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#759 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#759 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#760 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#760 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0be, 10'h000, 12'h30e, 12'hfff};
#760 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#761 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#761 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#762 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#762 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#763 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#763 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#764 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#764 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bf, 10'h000, 12'h30f, 12'hfff};
#764 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#765 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#765 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#765 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00b, 4'h3, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0bf, 10'h000, 12'h30f, 12'hfff};
#766 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#766 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#767 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#767 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#768 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#768 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c0, 10'h000, 12'h000, 12'hf00};
#768 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#769 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#769 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#769 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c0, 10'h000, 12'h000, 12'hf00};
#770 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#770 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#771 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001a0, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h000001a0, 5'h09, 32'h000001a0, 32'h00004940, 32'h00000005, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#771 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001a0, 32'h00000000, 32'h0000000d};
#772 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000068, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000068, 5'h0a, 32'h00000068, 32'h000050c0, 32'h00000003, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#772 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c1, 10'h000, 12'h001, 12'hf00};
#772 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000068, 32'h00000000, 32'h0000000d};
#773 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000208, 1'b0, 32'h00000000, 32'h00000068, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001a0, 32'h00000068, 32'h00000208, 5'h09, 32'h00000208, 32'h00004820, 32'h000001a0, 32'h00000068, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#773 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000208, 32'h00000000, 32'h00000068};
#774 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000215, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000208, 32'h0000000d, 32'h00000215, 5'h09, 32'h00000215, 32'h00004820, 32'h00000208, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#774 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000215, 32'h00000000, 32'h0000000d};
#775 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000854, 1'b0, 32'h00000000, 32'h00000215, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000215, 32'h00000854, 5'h09, 32'h00000854, 32'h00004880, 32'h00000002, 32'h00000215, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#775 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000854, 32'h00000000, 32'h00000215};
#776 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020854, 1'b0, 32'h00000002, 32'h00000854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000854, 32'h10020854, 5'h08, 32'h10020854, 32'h00004020, 32'h10020000, 32'h00000854, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#776 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020854, 32'h00000002, 32'h00000854};
#776 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c2, 10'h000, 12'h002, 12'hf00};
#777 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020854, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020854, 32'h00000003, 32'h10020854, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020854, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#777 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020854, 32'h00000002, 32'h00000003};
#777 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c2, 10'h000, 12'h002, 12'hf00};
#778 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#778 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#778 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c2, 10'h000, 12'h002, 12'hf00};
#779 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020854, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#779 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020854};
#780 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000854, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000854, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#780 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000854};
#780 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c3, 10'h000, 12'h003, 12'hf00};
#781 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000068, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000068, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#781 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000068};
#782 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#782 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#783 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#783 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#784 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000e, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000d, 32'h0000000d, 32'h0000000e, 5'h05, 32'h0000000e, 32'h00000001, 32'h0000000d, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#784 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c4, 10'h000, 12'h004, 12'hf00};
#784 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000e, 32'h00000000, 32'h0000000d};
#785 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000e, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000d, 32'h0000000d, 32'h0000000e, 5'h06, 32'h0000000e, 32'h00000001, 32'h0000000d, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#786 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000e, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000e, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#786 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#787 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#787 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#788 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#788 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c5, 10'h000, 12'h005, 12'hf00};
#788 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#789 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#789 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#790 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#790 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#791 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#791 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#791 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c5, 10'h000, 12'h005, 12'hf00};
#792 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#792 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#792 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c6, 10'h000, 12'h006, 12'hf00};
#793 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#793 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#794 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#794 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#795 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#795 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#795 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c6, 10'h000, 12'h006, 12'hf00};
#796 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#796 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c7, 10'h000, 12'h007, 12'hf00};
#796 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#797 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001c0, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h000001c0, 5'h09, 32'h000001c0, 32'h00004940, 32'h00000005, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#797 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001c0, 32'h00000000, 32'h0000000e};
#798 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000070, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000070, 5'h0a, 32'h00000070, 32'h000050c0, 32'h00000003, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#798 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000070, 32'h00000000, 32'h0000000e};
#799 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000230, 1'b0, 32'h00000000, 32'h00000070, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001c0, 32'h00000070, 32'h00000230, 5'h09, 32'h00000230, 32'h00004820, 32'h000001c0, 32'h00000070, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#799 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000230, 32'h00000000, 32'h00000070};
#800 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000023e, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000230, 32'h0000000e, 32'h0000023e, 5'h09, 32'h0000023e, 32'h00004820, 32'h00000230, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#800 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000023e, 32'h00000000, 32'h0000000e};
#800 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c8, 10'h000, 12'h008, 12'hf00};
#801 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000008f8, 1'b0, 32'h00000000, 32'h0000023e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000023e, 32'h000008f8, 5'h09, 32'h000008f8, 32'h00004880, 32'h00000002, 32'h0000023e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#801 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000008f8, 32'h00000000, 32'h0000023e};
#802 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100208f8, 1'b0, 32'h00000003, 32'h000008f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000008f8, 32'h100208f8, 5'h08, 32'h100208f8, 32'h00004020, 32'h10020000, 32'h000008f8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#802 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100208f8, 32'h00000003, 32'h000008f8};
#803 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100208f8, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100208f8, 32'h00000002, 32'h100208f8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100208f8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#803 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100208f8, 32'h00000003, 32'h00000002};
#803 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c8, 10'h000, 12'h008, 12'hf00};
#804 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#804 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#804 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0c9, 10'h000, 12'h009, 12'hf00};
#805 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100208f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100208f8, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#805 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100208f8};
#806 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000008f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000008f8, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#806 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000008f8};
#807 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000070, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000070, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#807 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000070};
#808 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#808 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#808 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ca, 10'h000, 12'h00a, 12'hf00};
#809 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#809 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#810 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#810 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#811 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#811 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#812 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#812 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cb, 10'h000, 12'h00b, 12'hf00};
#812 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#813 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#813 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#814 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#814 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#815 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#815 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#815 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cb, 10'h000, 12'h00b, 12'hf00};
#816 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#816 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#816 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cc, 10'h000, 12'h00c, 12'hf00};
#817 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#817 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#818 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#818 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#819 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#819 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#819 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cc, 10'h000, 12'h00c, 12'hf00};
#820 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#820 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cd, 10'h000, 12'h00d, 12'hf00};
#820 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#821 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001c0, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h000001c0, 5'h09, 32'h000001c0, 32'h00004940, 32'h00000005, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#821 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001c0, 32'h00000000, 32'h0000000e};
#822 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000070, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000070, 5'h0a, 32'h00000070, 32'h000050c0, 32'h00000003, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#822 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000070, 32'h00000000, 32'h0000000e};
#823 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000230, 1'b0, 32'h00000000, 32'h00000070, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001c0, 32'h00000070, 32'h00000230, 5'h09, 32'h00000230, 32'h00004820, 32'h000001c0, 32'h00000070, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#823 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000230, 32'h00000000, 32'h00000070};
#824 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h0000023e, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000230, 32'h0000000e, 32'h0000023e, 5'h09, 32'h0000023e, 32'h00004820, 32'h00000230, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#824 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000023e, 32'h00000000, 32'h0000000e};
#824 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ce, 10'h000, 12'h00e, 12'hf00};
#825 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h000008f8, 1'b0, 32'h00000000, 32'h0000023e, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000023e, 32'h000008f8, 5'h09, 32'h000008f8, 32'h00004880, 32'h00000002, 32'h0000023e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#825 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000008f8, 32'h00000000, 32'h0000023e};
#826 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h100208f8, 1'b0, 32'h00000002, 32'h000008f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000008f8, 32'h100208f8, 5'h08, 32'h100208f8, 32'h00004020, 32'h10020000, 32'h000008f8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#826 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100208f8, 32'h00000002, 32'h000008f8};
#827 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h100208f8, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100208f8, 32'h00000003, 32'h100208f8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100208f8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#827 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h100208f8, 32'h00000002, 32'h00000003};
#827 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ce, 10'h000, 12'h00e, 12'hf00};
#828 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#828 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#828 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00c, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0cf, 10'h000, 12'h00f, 12'hf00};
#829 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h100208f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100208f8, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#829 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h100208f8};
#830 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h000008f8, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000008f8, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#830 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h000008f8};
#831 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000070, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000070, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#831 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000070};
#832 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#832 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#832 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d0, 10'h000, 12'h000, 12'hf00};
#833 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#833 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#834 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h0000000f, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000e, 32'h0000000e, 32'h0000000f, 5'h05, 32'h0000000f, 32'h00000001, 32'h0000000e, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#834 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000000f, 32'h00000000, 32'h0000000e};
#835 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h0000000f, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000e, 32'h0000000e, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00000001, 32'h0000000e, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#836 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h0000000f, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h0000000f, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#836 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#836 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d1, 10'h000, 12'h001, 12'hf00};
#837 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#837 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#838 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#838 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#839 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#839 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#840 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#840 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d2, 10'h000, 12'h002, 12'hf00};
#840 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#841 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#841 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#841 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d2, 10'h000, 12'h002, 12'hf00};
#842 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#842 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#843 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#843 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#844 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#844 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d3, 10'h000, 12'h003, 12'hf00};
#844 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#845 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#845 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#845 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d3, 10'h000, 12'h003, 12'hf00};
#846 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#846 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#847 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001e0, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#847 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001e0, 32'h00000000, 32'h0000000f};
#848 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000078, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#848 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d4, 10'h000, 12'h004, 12'hf00};
#848 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000078, 32'h00000000, 32'h0000000f};
#849 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000258, 1'b0, 32'h00000000, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#849 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000258, 32'h00000000, 32'h00000078};
#850 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000267, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h0000000f, 32'h00000267, 5'h09, 32'h00000267, 32'h00004820, 32'h00000258, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#850 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000267, 32'h00000000, 32'h0000000f};
#851 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000099c, 1'b0, 32'h00000000, 32'h00000267, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000267, 32'h0000099c, 5'h09, 32'h0000099c, 32'h00004880, 32'h00000002, 32'h00000267, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#851 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000099c, 32'h00000000, 32'h00000267};
#852 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002099c, 1'b0, 32'h00000001, 32'h0000099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000099c, 32'h1002099c, 5'h08, 32'h1002099c, 32'h00004020, 32'h10020000, 32'h0000099c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#852 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002099c, 32'h00000001, 32'h0000099c};
#852 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d5, 10'h000, 12'h005, 12'hf00};
#853 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002099c, 1'b1, 32'h00000001, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002099c, 32'h00000002, 32'h1002099c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002099c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#853 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002099c, 32'h00000001, 32'h00000002};
#853 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d5, 10'h000, 12'h005, 12'hf00};
#854 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#854 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#854 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d5, 10'h000, 12'h005, 12'hf00};
#855 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002099c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#855 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002099c};
#856 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000099c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#856 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000099c};
#856 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d6, 10'h000, 12'h006, 12'hf00};
#857 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#857 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000078};
#858 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#858 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#859 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#859 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#860 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#860 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d7, 10'h000, 12'h007, 12'hf00};
#860 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#861 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#861 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#862 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#862 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#863 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#863 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#864 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#864 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d8, 10'h000, 12'h008, 12'hf00};
#864 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#865 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#865 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#865 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d8, 10'h000, 12'h008, 12'hf00};
#866 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#866 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#867 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#867 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#868 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#868 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d9, 10'h000, 12'h009, 12'hf00};
#868 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#869 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#869 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#869 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0d9, 10'h000, 12'h009, 12'hf00};
#870 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#870 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#871 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h000001e0, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#871 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000001e0, 32'h00000000, 32'h0000000f};
#872 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000078, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#872 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0da, 10'h000, 12'h00a, 12'hf00};
#872 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000078, 32'h00000000, 32'h0000000f};
#873 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000258, 1'b0, 32'h00000000, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#873 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000258, 32'h00000000, 32'h00000078};
#874 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000267, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h0000000f, 32'h00000267, 5'h09, 32'h00000267, 32'h00004820, 32'h00000258, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#874 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000267, 32'h00000000, 32'h0000000f};
#875 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h0000099c, 1'b0, 32'h00000000, 32'h00000267, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000267, 32'h0000099c, 5'h09, 32'h0000099c, 32'h00004880, 32'h00000002, 32'h00000267, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#875 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h0000099c, 32'h00000000, 32'h00000267};
#876 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h1002099c, 1'b0, 32'h00000002, 32'h0000099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h0000099c, 32'h1002099c, 5'h08, 32'h1002099c, 32'h00004020, 32'h10020000, 32'h0000099c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#876 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002099c, 32'h00000002, 32'h0000099c};
#876 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0db, 10'h000, 12'h00b, 12'hf00};
#877 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h1002099c, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h1002099c, 32'h00000003, 32'h1002099c, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h1002099c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#877 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h1002099c, 32'h00000002, 32'h00000003};
#877 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0db, 10'h000, 12'h00b, 12'hf00};
#878 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#878 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#878 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0db, 10'h000, 12'h00b, 12'hf00};
#879 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h1002099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h1002099c, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#879 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h1002099c};
#880 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h0000099c, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000099c, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#880 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h0000099c};
#880 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0dc, 10'h000, 12'h00c, 12'hf00};
#881 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#881 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000078};
#882 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#882 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#883 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#883 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#884 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000f, 32'h0000000f, 32'h00000010, 5'h05, 32'h00000010, 32'h00000001, 32'h0000000f, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#884 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0dd, 10'h000, 12'h00d, 12'hf00};
#884 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000010, 32'h00000000, 32'h0000000f};
#885 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h0000000f, 32'h0000000f, 32'h00000010, 5'h06, 32'h00000010, 32'h00000001, 32'h0000000f, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#886 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000010, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000010, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#886 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#887 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#887 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#888 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#888 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0de, 10'h000, 12'h00e, 12'hf00};
#888 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#889 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#889 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#890 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#890 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#891 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#891 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#891 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0de, 10'h000, 12'h00e, 12'hf00};
#892 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#892 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#892 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0df, 10'h000, 12'h00f, 12'hf00};
#893 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#893 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#894 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#894 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#895 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#895 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#895 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00d, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0df, 10'h000, 12'h00f, 12'hf00};
#896 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#896 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e0, 10'h000, 12'h000, 12'hf00};
#896 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#897 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000200, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000200, 5'h09, 32'h00000200, 32'h00004940, 32'h00000005, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#897 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000200, 32'h00000000, 32'h00000010};
#898 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000080, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000080, 5'h0a, 32'h00000080, 32'h000050c0, 32'h00000003, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#898 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000080, 32'h00000000, 32'h00000010};
#899 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000280, 1'b0, 32'h00000000, 32'h00000080, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000200, 32'h00000080, 32'h00000280, 5'h09, 32'h00000280, 32'h00004820, 32'h00000200, 32'h00000080, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#899 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000280, 32'h00000000, 32'h00000080};
#900 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000290, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000280, 32'h00000010, 32'h00000290, 5'h09, 32'h00000290, 32'h00004820, 32'h00000280, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#900 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000290, 32'h00000000, 32'h00000010};
#900 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e1, 10'h000, 12'h001, 12'hf00};
#901 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000a40, 1'b0, 32'h00000000, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000290, 32'h00000a40, 5'h09, 32'h00000a40, 32'h00004880, 32'h00000002, 32'h00000290, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#901 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000a40, 32'h00000000, 32'h00000290};
#902 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020a40, 1'b0, 32'h00000002, 32'h00000a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000a40, 32'h10020a40, 5'h08, 32'h10020a40, 32'h00004020, 32'h10020000, 32'h00000a40, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#902 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020a40, 32'h00000002, 32'h00000a40};
#903 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020a40, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020a40, 32'h00000002, 32'h10020a40, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020a40, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#903 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020a40, 32'h00000002, 32'h00000002};
#903 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e1, 10'h000, 12'h001, 12'hf00};
#904 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#904 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e2, 10'h000, 12'h002, 12'hf00};
#904 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#905 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020a40, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#905 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020a40};
#906 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000a40, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#906 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000a40};
#907 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000080, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000080, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#907 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000080};
#908 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#908 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#908 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e3, 10'h000, 12'h003, 12'hf00};
#909 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#909 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#910 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#910 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#911 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#911 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#912 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#912 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e4, 10'h000, 12'h004, 12'hf00};
#912 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#913 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#913 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#914 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#914 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#915 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#915 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#915 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e4, 10'h000, 12'h004, 12'hf00};
#916 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#916 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#916 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e5, 10'h000, 12'h005, 12'hf00};
#917 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#917 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#918 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#918 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#919 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#919 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#919 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e5, 10'h000, 12'h005, 12'hf00};
#920 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#920 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e6, 10'h000, 12'h006, 12'hf00};
#920 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#921 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000200, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000200, 5'h09, 32'h00000200, 32'h00004940, 32'h00000005, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#921 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000200, 32'h00000000, 32'h00000010};
#922 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000080, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000080, 5'h0a, 32'h00000080, 32'h000050c0, 32'h00000003, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#922 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000080, 32'h00000000, 32'h00000010};
#923 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h00000280, 1'b0, 32'h00000000, 32'h00000080, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000200, 32'h00000080, 32'h00000280, 5'h09, 32'h00000280, 32'h00004820, 32'h00000200, 32'h00000080, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#923 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000280, 32'h00000000, 32'h00000080};
#924 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h00000290, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000280, 32'h00000010, 32'h00000290, 5'h09, 32'h00000290, 32'h00004820, 32'h00000280, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#924 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000290, 32'h00000000, 32'h00000010};
#924 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e7, 10'h000, 12'h007, 12'hf00};
#925 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000a40, 1'b0, 32'h00000000, 32'h00000290, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000290, 32'h00000a40, 5'h09, 32'h00000a40, 32'h00004880, 32'h00000002, 32'h00000290, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#925 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000a40, 32'h00000000, 32'h00000290};
#926 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020a40, 1'b0, 32'h00000002, 32'h00000a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000a40, 32'h10020a40, 5'h08, 32'h10020a40, 32'h00004020, 32'h10020000, 32'h00000a40, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#926 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020a40, 32'h00000002, 32'h00000a40};
#927 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020a40, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020a40, 32'h00000003, 32'h10020a40, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020a40, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#927 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020a40, 32'h00000002, 32'h00000003};
#927 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e7, 10'h000, 12'h007, 12'hf00};
#928 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#928 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#928 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e8, 10'h000, 12'h008, 12'hf00};
#929 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020a40, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#929 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020a40};
#930 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000a40, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000a40, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#930 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000a40};
#931 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000080, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000080, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#931 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000080};
#932 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#932 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#932 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0e9, 10'h000, 12'h009, 12'hf00};
#933 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#933 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#934 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000011, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000010, 32'h00000010, 32'h00000011, 5'h05, 32'h00000011, 32'h00000001, 32'h00000010, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#934 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000011, 32'h00000000, 32'h00000010};
#935 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000011, 1'b0, 32'h00000000, 32'h00000010, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000010, 32'h00000010, 32'h00000011, 5'h06, 32'h00000011, 32'h00000001, 32'h00000010, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#936 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000011, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000011, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#936 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#936 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ea, 10'h000, 12'h00a, 12'hf00};
#937 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#937 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#938 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#938 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#939 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#939 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#940 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#940 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0eb, 10'h000, 12'h00b, 12'hf00};
#940 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#941 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#941 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#941 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0eb, 10'h000, 12'h00b, 12'hf00};
#942 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#942 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#943 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#943 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#944 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#944 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ec, 10'h000, 12'h00c, 12'hf00};
#944 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#945 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#945 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#945 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ec, 10'h000, 12'h00c, 12'hf00};
#946 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#946 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#947 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000220, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000011, 32'h00000220, 5'h09, 32'h00000220, 32'h00004940, 32'h00000005, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#947 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000220, 32'h00000000, 32'h00000011};
#948 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000088, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000011, 32'h00000088, 5'h0a, 32'h00000088, 32'h000050c0, 32'h00000003, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#948 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ed, 10'h000, 12'h00d, 12'hf00};
#948 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000088, 32'h00000000, 32'h00000011};
#949 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000002a8, 1'b0, 32'h00000000, 32'h00000088, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000220, 32'h00000088, 32'h000002a8, 5'h09, 32'h000002a8, 32'h00004820, 32'h00000220, 32'h00000088, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#949 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000002a8, 32'h00000000, 32'h00000088};
#950 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000002b9, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000002a8, 32'h00000011, 32'h000002b9, 5'h09, 32'h000002b9, 32'h00004820, 32'h000002a8, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#950 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000002b9, 32'h00000000, 32'h00000011};
#951 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000ae4, 1'b0, 32'h00000000, 32'h000002b9, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000002b9, 32'h00000ae4, 5'h09, 32'h00000ae4, 32'h00004880, 32'h00000002, 32'h000002b9, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#951 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000ae4, 32'h00000000, 32'h000002b9};
#952 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020ae4, 1'b0, 32'h00000000, 32'h00000ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000ae4, 32'h10020ae4, 5'h08, 32'h10020ae4, 32'h00004020, 32'h10020000, 32'h00000ae4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#952 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020ae4, 32'h00000000, 32'h00000ae4};
#952 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ee, 10'h000, 12'h00e, 12'hf00};
#953 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020ae4, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020ae4, 32'h00000002, 32'h10020ae4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020ae4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#953 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020ae4, 32'h00000000, 32'h00000002};
#953 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ee, 10'h000, 12'h00e, 12'hf00};
#954 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000d0};
#954 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000d0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'h1f, 32'h004000d0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#954 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ee, 10'h000, 12'h00e, 12'hf00};
#955 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020ae4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#955 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020ae4};
#956 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000ae4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#956 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000ae4};
#956 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00e, 4'h0, 1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h0, 4'h0, 10'h0ef, 10'h000, 12'h00f, 12'hf00};
#957 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000088, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000088, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#957 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000088};
#958 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#958 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#959 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000d0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#959 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#960 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d0, 32'h24040032, 32'h00000032, 1'b0, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000032, 5'h04, 32'h00000032, 32'h00000032, 32'h00000000, 32'h00000032, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#960 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f0, 10'h000, 12'h100, 12'h0f0};
#960 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000032, 32'h00000000, 32'h00000002};
#961 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d4, 32'h00000000, 32'h00000000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h00, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#961 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
#962 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000d8, 32'h24040003, 32'h00000003, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000032, 32'h00000003, 5'h04, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#962 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000003, 32'h00000000, 32'h00000032};
#963 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000dc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000e0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#963 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#964 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#964 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f1, 10'h000, 12'h101, 12'h0f0};
#964 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#965 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000d0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#965 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000d0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000d0, 32'h004000e0};
#965 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f1, 10'h000, 12'h101, 12'h0f0};
#966 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#966 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#967 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#967 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#968 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#968 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f2, 10'h000, 12'h102, 12'h0f0};
#968 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#969 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#969 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#969 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f2, 10'h000, 12'h102, 12'h0f0};
#970 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#970 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#971 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000220, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000011, 32'h00000220, 5'h09, 32'h00000220, 32'h00004940, 32'h00000005, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#971 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000220, 32'h00000000, 32'h00000011};
#972 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000088, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000011, 32'h00000088, 5'h0a, 32'h00000088, 32'h000050c0, 32'h00000003, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#972 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f3, 10'h000, 12'h103, 12'h0f0};
#972 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000088, 32'h00000000, 32'h00000011};
#973 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000002a8, 1'b0, 32'h00000000, 32'h00000088, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000220, 32'h00000088, 32'h000002a8, 5'h09, 32'h000002a8, 32'h00004820, 32'h00000220, 32'h00000088, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#973 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000002a8, 32'h00000000, 32'h00000088};
#974 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h01254820, 32'h000002b9, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000002a8, 32'h00000011, 32'h000002b9, 5'h09, 32'h000002b9, 32'h00004820, 32'h000002a8, 32'h00000011, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#974 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000002b9, 32'h00000000, 32'h00000011};
#975 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'h00094880, 32'h00000ae4, 1'b0, 32'h00000000, 32'h000002b9, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000002b9, 32'h00000ae4, 5'h09, 32'h00000ae4, 32'h00004880, 32'h00000002, 32'h000002b9, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#975 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000ae4, 32'h00000000, 32'h000002b9};
#976 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'h01094020, 32'h10020ae4, 1'b0, 32'h00000002, 32'h00000ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000ae4, 32'h10020ae4, 5'h08, 32'h10020ae4, 32'h00004020, 32'h10020000, 32'h00000ae4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#976 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020ae4, 32'h00000002, 32'h00000ae4};
#976 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f4, 10'h000, 12'h104, 12'h0f0};
#977 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'had040000, 32'h10020ae4, 1'b1, 32'h00000002, 32'h00000003, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10020ae4, 32'h00000003, 32'h10020ae4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020ae4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#977 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h10020ae4, 32'h00000002, 32'h00000003};
#977 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f4, 10'h000, 12'h104, 12'h0f0};
#978 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000e0};
#978 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h004000e0, 32'h004000e0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000e0, 32'h10010ffc, 5'h1f, 32'h004000e0, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#978 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f4, 10'h000, 12'h104, 12'h0f0};
#979 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'h00000001, 32'h10020ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020ae4, 32'h10010ff8, 5'h08, 32'h00000001, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#979 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h10020ae4};
#980 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hffffffff, 32'h00000ae4, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000ae4, 32'h10010ff4, 5'h09, 32'hffffffff, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#980 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'h00000ae4};
#980 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f5, 10'h000, 12'h105, 12'h0f0};
#981 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'h00000004, 32'h00000088, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000088, 32'h10010ff0, 5'h0a, 32'h00000004, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#981 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000088};
#982 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000009, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#982 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000009, 32'h10010ff0};
#983 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h004000e0, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'h0000000X, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#983 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#984 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e0, 32'h20a50001, 32'h00000012, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000011, 32'h00000011, 32'h00000012, 5'h05, 32'h00000012, 32'h00000001, 32'h00000011, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#984 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f6, 10'h000, 12'h106, 12'h0f0};
#984 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000012, 32'h00000000, 32'h00000011};
#985 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e4, 32'h20c60001, 32'h00000012, 1'b0, 32'h00000000, 32'h00000011, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000011, 32'h00000011, 32'h00000012, 5'h06, 32'h00000012, 32'h00000001, 32'h00000011, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#986 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000e8, 32'h28c8001e, 32'h00000001, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'b1x011, 1'b0, 32'h00000012, 32'h00000001, 32'h00000001, 5'h08, 32'h00000001, 32'h0000001e, 32'h00000012, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#986 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000001};
#987 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ec, 32'h1500fff6, 32'h00000001, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff6, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#987 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000};
#988 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000c8, 32'h24040002, 32'h00000002, 1'b0, 32'h00000000, 32'h00000003, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#988 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f7, 10'h000, 12'h107, 12'h0f0};
#988 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h00000002, 32'h00000000, 32'h00000003};
#989 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000cc, 32'h0c10005c, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00400104, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00400104, 32'hxxxxxxxx, 5'h1f, 32'h004000d0, 32'h0000005c, 32'hxxxxxxxx, 32'h00X00XXX, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#989 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h0000000X, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00400104};
#990 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400170, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000004, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#990 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h10011000};
#991 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400174, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h004000e0, 32'h004000d0, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h004000d0, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#991 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h004000e0, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h004000e0, 32'h004000d0};
#991 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f7, 10'h000, 12'h107, 12'h0f0};
#992 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000001, 32'h00000001};
#992 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400178, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000001, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#992 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f8, 10'h000, 12'h108, 12'h0f0};
#993 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040017c, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hffffffff, 32'hffffffff, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hffffffff, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#993 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hffffffff, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'hffffffff, 32'hffffffff};
#994 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400180, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000004, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#994 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000004, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000004, 32'h00000004};
#995 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400184, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000003, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#995 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h10020000};
#995 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f8, 10'h000, 12'h108, 12'h0f0};
#996 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400188, 32'h34280000, 32'h10020000, 1'b0, 32'h00000003, 32'h00000001, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'h00000001, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#996 {smem_addr, charcode, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_addr, bmem_color} <= {11'h00f, 4'h1, 1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0f9, 10'h000, 12'h109, 12'h0f0};
#996 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000009, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000003, 32'h00000001};
#997 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040018c, 32'h00064940, 32'h00000240, 1'b0, 32'h00000000, 32'h00000012, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000012, 32'h00000240, 5'h09, 32'h00000240, 32'h00004940, 32'h00000005, 32'h00000012, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#997 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000240, 32'h00000000, 32'h00000012};
#998 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400190, 32'h000650c0, 32'h00000090, 1'b0, 32'h00000000, 32'h00000012, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000012, 32'h00000090, 5'h0a, 32'h00000090, 32'h000050c0, 32'h00000003, 32'h00000012, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#998 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h00000090, 32'h00000000, 32'h00000012};
#999 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400194, 32'h012a4820, 32'h000002d0, 1'b0, 32'h00000000, 32'h00000090, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000240, 32'h00000090, 32'h000002d0, 5'h09, 32'h000002d0, 32'h00004820, 32'h00000240, 32'h00000090, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#999 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'h000002d0, 32'h00000000, 32'h00000090};

join
end

endmodule